`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/13/2022 11:21:25 PM
// Design Name: 
// Module Name: TB
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TB_new();
reg clk_100=0;
reg clk_166=0;
reg [7:0]r=0,g=0,b=0;
reg wr_en;
reg reset=0,start_kmeans=0;
reg start_lab_conv=0;
wire [2:0]EB_LB_HD;
wire NN_done;

wire done_features;
wire finish_lab,done_kmeans;
wire HS,VS,done,done_cluster_settings;
wire [3:0]blue,green,red;
 
 design_sim_wrapper uut
   (EB_LB_HD,
  NN_done,
  b,
  clk_100,
  done,
  done_cluster_settings,
  done_features,
  done_kmeans,
  finish_lab,
  g,
  r,
  reset,
  wr_en);

int R[2500]; 
int G[2500]; 
int B[2500];
int i = 0;
initial begin
/*
  R = '{181,  170,  169,  165,  162,  147,  153,  159,  150,  141,
  158,  108,  156,  155,  158,  120,   60,  122,  161,  149,
  176,  137,  143,  150,  161,  132,   89,  100,  121,  158,
  193,  165,  145,  125,  157,  135,  120,  112,   87,  155,
  198,  166,  164,  116,  136,  148,  130,  114,   97,  146,
  201,  165,  166,  157,  130,  149,  129,  106,   94,  113,
  204,  189,  163,  164,  140,  133,  120,   98,   68,  100,
  202,  197,  169,  156,  147,  135,  120,   89,   65,  137,
  200,  200,  192,  168,  140,  120,  121,  104,   60,  121,
  199,  197,  196,  195,  187,  166,  160,  161,  153,  137};

  G = '{
  175,  162,  163,  160,  155,  139,  143,  150,  142,  133,
  147,  101,  167,  168,  166,  130,   66,  116,  150,  139,
  170,  137,  158,  167,  171,  130,  104,  114,  112,  146,
  188,  176,  161,  147,  163,  125,  135,  137,   86,  143,
  191,  173,  177,  131,  153,  154,  139,  138,  106,  134,
  193,  166,  181,  151,  135,  154,  145,  128,  115,  104,
  197,  186,  174,  156,  125,  148,  137,  102,   76,   91,
  195,  189,  175,  173,  164,  154,  139,  102,   64,  125,
  193,  190,  184,  173,  157,  143,  143,  127,   64,  114,
  193,  190,  187,  183,  179,  165,  157,  156,  145,  130};

  B = '{181,  166,  159,  153,  151,  143,  152,  157,  149,  140,
  142,   60,  120,  124,  121,   86,   42,  115,  157,  145,
  160,   92,  118,  128,  135,   94,   56,   72,  111,  153,
  184,  131,  123,  104,  133,   97,   88,   83,   65,  149,
  192,  134,  142,   90,  107,  115,   97,   85,   67,  137,
  198,  142,  145,  128,   94,  106,   96,   77,   66,  102,
  201,  172,  134,  131,   99,   96,   79,   63,   38,   91,
  197,  190,  145,  134,  123,  110,   91,   53,   37,  128,
  195,  194,  183,  148,  117,   98,   96,   82,   35,  103,
  196,  193,  192,  189,  176,  150,  142,  146,  136,  116};
*/
R = '{
182, 178, 184, 180, 178, 175, 177, 179, 177, 177, 171, 173, 173, 170, 173, 174, 171, 172, 171, 166, 167, 169, 174, 166, 167, 167, 172, 162, 152, 152, 162, 168, 169, 156, 148, 154, 152, 163, 156, 145, 154, 151, 147, 152, 146, 141, 135, 134, 141, 136,  
   185, 186, 185, 178, 180, 175, 176, 177, 175, 177, 176, 174, 171, 168, 173, 171, 168, 170, 171, 164, 168, 166, 174, 160, 168, 167, 164, 158, 158, 156, 155, 163, 165, 161, 155, 156, 155, 159, 156, 149, 148, 148, 145, 147, 147, 144, 138, 139, 139, 143,  
   186, 187, 183, 179, 178, 177, 175, 178, 178, 178, 180, 176, 170, 173, 174, 166, 163, 172, 169, 163, 168, 169, 172, 164, 170, 172, 171, 171, 156, 159, 157, 162, 158, 160, 159, 154, 158, 156, 161, 154, 154, 152, 150, 146, 145, 152, 144, 142, 137, 136,  
   190, 184, 179, 181, 181, 185, 183, 181, 179, 176, 176, 175, 175, 177, 175, 172, 168, 169, 177, 171, 169, 159, 157, 164, 159, 175, 162, 169, 170, 163, 162, 161, 159, 158, 156, 162, 158, 155, 155, 158, 159, 155, 154, 151, 144, 147, 147, 145, 144, 136,  
   189, 185, 184, 184, 170, 167, 177, 182, 171, 168, 168, 159, 147, 141, 136, 147, 141, 134, 149, 153, 160, 155, 144, 127,  89,  72,  76,  98, 101, 114, 139, 159, 164, 161, 160, 166, 167, 161, 151, 156, 161, 161, 153, 149, 144, 145, 144, 146, 145, 143,  
   184, 183, 186, 175, 101,  78,  81,  87,  51,  92, 155, 154, 156, 146, 130, 136, 136, 140, 136, 152, 157, 156, 166, 162, 151, 137,  98,  49,  27,  34,  41,  51,  63,  97, 145, 165, 163, 156, 157, 153, 155, 164, 159, 152, 147, 142, 146, 150, 145, 146,  
   184, 184, 189, 135,  66,  61,  84,  81,  97, 102, 166, 172, 166, 165, 156, 163, 161, 158, 154, 173, 157, 151, 167, 167, 152, 147, 152, 149,  96,  45,  33,  28,  31,  28,  45, 108, 155, 164, 160, 155, 162, 162, 160, 154, 148, 148, 148, 146, 151, 149,  
   185, 190, 191, 131,  80,  55,  87, 128, 164, 162, 155, 172, 159, 157, 170, 160, 156, 143, 159, 166, 139, 142, 170, 174, 158, 141, 151, 149, 151, 119,  62,  40,  41,  33,  24,  26,  69, 156, 166, 162, 170, 169, 159, 152, 149, 151, 148, 149, 152, 148,  
   184, 182, 191, 159,  61,  57,  49, 108, 153, 172, 155, 162, 136, 142, 162, 167, 151, 162, 174, 156, 151, 155, 143, 159, 175, 155, 164, 150, 142, 112,  48,  50,  56,  66,  58,  35,  22, 121, 169, 163, 168, 165, 156, 158, 156, 150, 148, 152, 152, 149,  
   182, 181, 185, 173,  85,  84,  72,  84, 139, 164, 157, 155, 158, 136, 149, 161, 155, 150, 168, 147, 169, 172, 154, 144, 170, 171, 159, 154, 143,  91,  31,  42,  42,  86,  93, 115,  63,  34,  92, 153, 163, 165, 160, 158, 158, 156, 149, 150, 154, 153,  
   192, 188, 190, 173, 105, 106, 115, 125, 132, 156, 156, 151, 140, 139, 164, 156, 160, 142, 154, 148, 170, 168, 165, 148, 142, 146, 155, 156, 136,  76,  32,  41,  49,  90, 103, 128, 125,  60,  18,  72, 155, 163, 160, 152, 154, 154, 155, 153, 153, 150,  
   191, 191, 191, 181, 118,  89,  93, 117, 144, 166, 138, 148, 153, 142, 141, 159, 153, 156, 165, 158, 163, 160, 155, 164, 158, 167, 159, 159, 126,  70,  49,  49,  86, 121, 116, 108, 120, 130,  47,  22,  89, 166, 160, 155, 158, 158, 156, 155, 154, 149,  
   193, 191, 192, 189, 131, 116, 133, 136, 135, 164, 140, 135, 153, 140, 125, 144, 152, 165, 153, 165, 162, 153, 163, 168, 164, 156, 153, 174, 135,  51,  40,  72, 113, 114, 121, 129, 129, 140, 107,  27,  27, 104, 157, 158, 157, 158, 155, 153, 155, 154,  
   194, 194, 196, 193, 147, 149, 138, 142, 171, 169, 163, 111, 110, 138, 135, 130, 144, 148, 142, 157, 153, 156, 154, 161, 141, 146, 155, 156, 120,  74,  39,  92, 131, 110, 120, 133, 131, 136, 137,  61,  24,  31, 123, 164, 153, 157, 153, 156, 153, 152,  
   193, 192, 194, 197, 150, 146, 150, 153, 170, 166, 162, 136,  98, 138, 164, 141, 127, 131, 128, 137, 158, 154, 157, 158, 165, 129, 159, 155, 117,  90,  68,  94, 124, 111, 115, 121, 124, 136, 139, 116,  30,  23,  67, 158, 153, 156, 157, 159, 152, 149,  
   197, 194, 192, 199, 167, 133, 154, 168, 162, 158, 164, 166, 130, 105, 142, 149, 130, 131, 132, 135, 153, 157, 164, 162, 175, 151, 157, 171, 148,  91, 100, 114, 124, 122, 104,  98, 110, 123, 129, 140,  61,  23,  34, 136, 156, 154, 153, 156, 154, 151,  
   199, 197, 196, 201, 179, 127, 145, 162, 171, 177, 169, 161, 145, 102, 107, 164, 154, 136, 130, 140, 150, 157, 147, 153, 171, 150, 149, 159, 101, 106, 135, 129, 111, 136, 101,  93, 113, 120, 125, 127, 109,  27,  23,  97, 167, 159, 161, 159, 156, 153,  
   198, 200, 202, 207, 190, 141, 145, 160, 172, 169, 168, 162, 158, 125,  81, 105, 146, 161, 139, 118, 141, 157, 152, 151, 165, 162, 135, 138, 102, 112, 127, 146, 111, 120,  98,  93, 100, 122, 125, 113, 136,  52,  25,  55, 158, 162, 160, 155, 153, 155,  
   197, 197, 204, 206, 191, 149, 153, 159, 173, 172, 165, 166, 139, 142, 110,  89,  97, 139, 150, 144, 145, 151, 154, 167, 177, 163, 137, 107, 113, 118, 139, 164, 139, 118, 123,  89,  94, 112, 118, 116, 145, 100,  28,  29, 125, 159, 157, 153, 154, 153,  
   198, 199, 202, 202, 197, 157, 152, 154, 169, 168, 181, 179, 165, 157, 135,  97,  91,  88, 118, 156, 145, 150, 156, 167, 172, 158, 144, 115, 107, 120, 146, 138, 129, 135, 125, 106,  99, 117, 116, 113, 134, 125,  32,  24, 107, 164, 155, 158, 160, 154,  
   199, 200, 200, 199, 200, 164, 152, 155, 168, 179, 175, 166, 173, 179, 144, 112, 104,  79,  75, 114, 144, 167, 151, 149, 151, 153, 156, 121, 106, 127, 143, 135, 121, 109, 121, 112, 104, 104, 106, 119, 117, 129,  46,  19,  93, 167, 160, 162, 154, 157,  
   200, 200, 203, 202, 201, 169, 146, 170, 172, 175, 177, 175, 162, 164, 154, 137, 133,  98,  94,  79, 126, 163, 149, 133, 146, 146, 147, 137, 116, 129, 125, 139, 142, 110, 114, 112, 104, 102, 116, 110, 111, 124,  91,  27,  90, 163, 159, 158, 156, 156,  
   201, 201, 199, 200, 204, 176, 151, 173, 170, 166, 167, 165, 173, 154, 165, 144, 110, 100,  96,  80,  89, 136, 170, 133, 145, 152, 146, 146, 142, 124, 139, 143, 130, 121, 119, 113, 100, 105, 123, 116, 106, 115, 128,  84,  37, 146, 164, 159, 159, 155,  
   201, 202, 198, 197, 201, 185, 147, 161, 168, 169, 170, 168, 148, 142, 167, 152, 128,  98, 108, 104,  97,  83, 141, 164, 149, 153, 144, 146, 158, 148, 151, 152, 141, 125, 116, 108, 122, 130, 117, 112,  97, 108, 125, 109,  24, 103, 169, 158, 160, 161,  
   200, 200, 199, 197, 197, 182, 136, 151, 164, 163, 177, 164, 175, 169, 167, 158, 147, 136, 133, 127, 121, 115, 118, 159, 162, 162, 147, 156, 183, 170, 147, 123, 128, 135, 109, 116, 123, 126, 137, 113,  93, 109, 131, 122,  36,  54, 158, 159, 157, 159,  
   200, 199, 196, 196, 198, 187,  92, 137, 160, 165, 168, 168, 158, 152, 192, 192, 157, 142, 123, 137, 116, 105, 126, 121, 149, 159, 155, 166, 189, 170, 156, 147, 123, 110, 103,  88, 116, 128, 127, 108,  92, 115, 124, 117,  44,  29, 134, 158, 157, 154,  
   201, 197, 199, 198, 197, 203, 115, 102, 182, 159, 153, 166, 167, 156, 169, 177, 168, 158, 147, 144, 118, 131, 129, 133, 129, 144, 163, 169, 174, 169, 159, 136, 137, 124, 103,  81,  97, 117, 121, 102, 111, 111, 114, 127,  47,  19,  88, 158, 161, 160,  
   200, 201, 199, 199, 199, 203, 154,  97, 171, 154, 158, 176, 164, 162, 172, 174, 169, 150, 174, 132, 117, 131, 135, 129, 133, 114, 126, 172, 155, 152, 139, 133, 126, 129, 103,  71,  96, 116, 126, 103, 106, 109, 119, 121,  45,  17,  54, 151, 157, 156,  
   205, 202, 200, 204, 203, 204, 194, 137, 168, 161, 158, 177, 180, 167, 169, 164, 156, 174, 170, 129, 119, 120, 130, 122, 152, 142, 103, 132, 157, 145, 130, 139, 136, 112, 105,  62,  76, 124, 128, 101, 111, 119, 112, 111,  42,  20,  31, 130, 157, 157,  
   202, 201, 202, 208, 207, 205, 208, 183, 165, 162, 168, 163, 172, 161, 160, 164, 170, 178, 184, 159, 161, 151, 146, 150, 150, 137, 126, 108, 131, 140, 135, 151, 146, 120, 105,  79,  76, 105, 120, 105, 116, 113, 108, 109,  37,  21,  23, 108, 157, 158,  
   205, 205, 196, 205, 206, 206, 204, 200, 155, 161, 177, 152, 155, 154, 168, 170, 171, 179, 165, 158,  98, 109, 163, 159, 148, 136, 126, 130, 112, 130, 136, 143, 152, 119, 112, 107, 124,  55,  80, 104, 108, 110, 115, 100,  27,  22,  20,  95, 160, 154,  
   206, 204, 200, 196, 198, 207, 200, 202, 178, 159, 165, 177, 163, 152, 154, 175, 198, 180, 152, 145, 108,  74, 122, 148, 157, 141, 133, 126, 125,  97, 117, 135, 148, 125, 108, 112, 142,  88,  76, 101,  86, 102, 116,  65,  18,  21,  21, 103, 164, 159,  
   206, 203, 201, 201, 198, 201, 201, 200, 185, 145, 160, 184, 176, 173, 161, 151, 172, 169, 162, 162, 184, 109, 113, 141, 156, 140, 137, 142, 130, 125,  95, 127, 142, 131, 125, 122, 148,  55,  25,  84, 110, 106, 112,  31,  15,  19,  24, 125, 162, 162,  
   202, 203, 203, 202, 197, 200, 199, 194, 194, 146, 158, 170, 172, 171, 143, 170, 165, 150, 152, 167, 164, 130, 112, 136, 148, 144, 149, 147, 146, 129, 105,  80, 100, 141, 134, 123, 150,  81,  11,  56, 119, 129, 112,  18,  16,  19,  30, 136, 158, 153,  
   202, 201, 199, 199, 202, 198, 198, 196, 197, 181, 141, 159, 162, 154, 163, 165, 158, 152, 163, 186, 163, 169, 138, 121, 122, 119, 142, 144, 147, 137, 134, 107,  59,  78, 131, 112, 129, 121,  19,  48, 117, 130,  95,  22,  18,  17,  60, 154, 153, 156,  
   204, 201, 201, 201, 201, 199, 199, 200, 198, 199, 155, 160, 167, 163, 166, 169, 159, 156, 162, 166, 164, 163, 157, 151, 147, 126, 144, 135, 132, 128, 143, 150, 109,  56,  62, 121, 113, 134,  93,  56,  91, 113,  66,  25,  20,  20, 109, 161, 154, 160,  
   203, 206, 202, 203, 197, 198, 200, 201, 201, 199, 178, 145, 173, 177, 162, 150, 153, 162, 168, 137, 161, 138, 153, 169, 153, 141, 135, 129, 123, 124, 132, 138, 136,  97,  48,  53, 110, 112, 123,  90,  95, 118,  38,  27,  20,  33, 144, 157, 157, 157,  
   199, 201, 202, 201, 201, 202, 199, 198, 195, 197, 195, 155, 146, 164, 164, 153, 158, 170, 154, 154, 151, 141, 158, 159, 158, 149, 134, 131, 125, 122, 131, 131, 130, 140, 102,  43,  43,  97, 108, 105,  99, 120,  64,  27,  19,  61, 157, 159, 162, 154,  
   200, 202, 203, 204, 206, 203, 198, 194, 191, 195, 196, 188, 159, 172, 175, 154, 158, 161, 156, 163, 150, 139, 137, 134, 152, 146, 146, 131, 119, 122, 137, 146, 141, 135, 140, 107,  56,  36,  66,  72,  99, 106,  98,  31,  22, 111, 161, 159, 159, 153,  
   198, 203, 199, 201, 202, 202, 196, 198, 193, 194, 197, 195, 189, 147, 151, 162, 163, 167, 158, 159, 144, 138, 134, 139, 154, 150, 136, 136, 129, 120, 120, 124, 132, 138, 128, 123, 110,  68,  37,  40,  57,  73,  98,  75, 122, 155, 155, 156, 157, 155,  
   199, 201, 199, 200, 203, 202, 201, 196, 195, 194, 194, 198, 194, 165, 135, 158, 154, 150, 141, 138, 125, 122, 138, 133, 138, 129, 119, 124, 118, 112, 123, 104, 135, 150, 144, 145, 143, 116,  87,  52,  29,  28,  22,  41, 135, 164, 160, 159, 156, 159,  
   199, 198, 197, 203, 204, 201, 201, 201, 198, 192, 195, 194, 200, 196, 177, 165, 155, 135, 145, 142, 137, 135, 137, 141, 133, 124, 128, 145, 122, 115, 120, 105, 131, 147, 149, 144, 127, 117, 126,  94,  46,  30,  28,  12,  30, 104, 156, 161, 158, 156,  
   200, 197, 199, 205, 203, 205, 203, 204, 200, 197, 202, 195, 189, 194, 198, 185, 174, 159, 159, 150, 164, 150, 138, 132, 127, 128, 122, 135, 105, 121, 101, 103, 123, 129, 120, 112,  92, 104, 117, 121,  85,  42,  40,  27,  12,  17, 107, 164, 166, 164,  
   201, 201, 200, 203, 208, 203, 198, 199, 197, 201, 198, 198, 195, 193, 203, 205, 198, 184, 160, 160, 133, 160, 141, 121, 116, 129, 128, 112, 113, 121,  99, 140, 124, 111, 105,  98, 103, 111, 106, 108, 112,  80,  56,  49,  20,  19, 111, 158, 110, 101,  
   199, 197, 196, 198, 202, 201, 195, 191, 199, 203, 200, 202, 197, 195, 195, 195, 194, 195, 189, 186, 159, 167, 146, 123, 120, 135, 121, 115, 122, 112, 119, 133, 114, 111, 124, 103, 108, 113, 102,  96, 100,  46,  37,  95,  76,  38, 121, 144,  80,  20,  
   199, 196, 201, 202, 195, 196, 194, 191, 195, 197, 197, 191, 192, 199, 192, 186, 194, 192, 195, 194, 193, 183, 172, 148, 137, 132, 127, 115, 107, 120, 117, 106,  99, 107, 126, 120, 111, 106, 101,  98,  86,  68,  91, 161, 157,  87, 120, 140,  76,  42,  
   200, 200, 199, 200, 198, 202, 204, 198, 195, 197, 197, 196, 200, 196, 194, 198, 198, 194, 195, 188, 187, 199, 198, 180, 182, 173, 152, 129, 129, 128, 116, 121, 129, 157, 170, 160, 152, 158, 161, 164, 166, 171, 171, 167, 178, 116, 103, 148, 123, 140,  
   198, 201, 201, 199, 196, 199, 195, 196, 199, 198, 198, 195, 199, 197, 194, 194, 194, 192, 195, 190, 188, 196, 197, 193, 194, 191, 192, 186, 183, 178, 178, 179, 184, 177, 178, 178, 173, 177, 174, 173, 172, 170, 161, 160, 171, 157, 135, 160, 164, 156,  
   200, 198, 200, 200, 198, 197, 195, 196, 198, 193, 193, 200, 198, 192, 190, 188, 193, 192, 198, 196, 192, 193, 196, 192, 196, 196, 191, 193, 189, 185, 184, 184, 180, 181, 179, 176, 175, 179, 176, 178, 176, 164, 161, 161, 161, 164, 160, 159, 157, 150,  
   203, 199, 198, 194, 197, 201, 198, 195, 188, 194, 195, 194, 201, 192, 194, 186, 189, 195, 198, 198, 194, 198, 193, 192, 188, 191, 189, 184, 185, 183, 187, 183, 179, 180, 184, 185, 178, 173, 174, 174, 174, 170, 161, 162, 164, 163, 160, 155, 152, 148  
};

G = '{
177, 173, 179, 175, 173, 170, 171, 172, 170, 170, 164, 166, 166, 163, 166, 167, 164, 165, 164, 160, 161, 162, 163, 155, 156, 156, 161, 151, 144, 146, 155, 158, 158, 144, 139, 147, 145, 156, 149, 138, 147, 144, 140, 145, 139, 134, 128, 127, 134, 129,
   180, 181, 180, 173, 175, 171, 170, 170, 168, 170, 169, 167, 164, 161, 166, 164, 161, 163, 164, 158, 162, 159, 163, 149, 157, 156, 154, 147, 151, 149, 148, 153, 154, 150, 146, 150, 148, 152, 149, 142, 141, 141, 138, 140, 140, 137, 131, 132, 132, 136,
   181, 182, 178, 174, 173, 171, 169, 171, 171, 171, 174, 169, 163, 165, 167, 159, 156, 166, 163, 157, 163, 163, 162, 153, 159, 161, 160, 160, 148, 152, 150, 153, 148, 150, 150, 147, 151, 149, 154, 147, 146, 145, 143, 139, 138, 145, 137, 135, 130, 129,
   183, 177, 172, 173, 173, 176, 176, 175, 171, 167, 168, 166, 167, 169, 165, 161, 157, 159, 166, 159, 158, 148, 148, 155, 149, 165, 151, 160, 160, 153, 152, 152, 151, 149, 146, 151, 148, 144, 144, 148, 149, 144, 144, 141, 137, 140, 140, 135, 133, 126,
   182, 177, 177, 178, 159, 149, 162, 169, 161, 157, 161, 158, 152, 150, 147, 157, 145, 129, 143, 155, 159, 151, 140, 122,  82,  69,  73,  94,  96, 108, 133, 149, 152, 149, 149, 155, 156, 150, 140, 145, 150, 150, 142, 139, 137, 138, 137, 135, 134, 132,
   177, 176, 179, 159,  72,  56,  65,  71,  42,  89, 157, 163, 167, 161, 152, 161, 157, 159, 154, 171, 171, 166, 177, 173, 162, 143, 100,  48,  26,  34,  40,  47,  58,  93, 137, 154, 152, 145, 146, 142, 144, 153, 148, 142, 140, 135, 138, 140, 134, 135,
   178, 177, 179, 113,  47,  53,  77,  74,  96, 106, 174, 182, 166, 164, 169, 177, 176, 176, 168, 182, 166, 165, 180, 177, 164, 162, 168, 157,  98,  45,  31,  28,  29,  27,  45, 103, 144, 152, 149, 144, 151, 151, 149, 143, 138, 139, 138, 135, 140, 138,
   180, 182, 180, 111,  67,  42,  77, 127, 167, 170, 164, 180, 160, 161, 184, 174, 172, 160, 172, 176, 147, 160, 187, 181, 153, 136, 164, 167, 164, 129,  70,  44,  36,  30,  25,  25,  63, 146, 155, 151, 159, 158, 148, 141, 138, 140, 137, 138, 141, 137,
   178, 174, 180, 140,  40,  40,  37, 106, 159, 183, 167, 173, 146, 156, 180, 182, 167, 179, 189, 169, 157, 164, 152, 170, 167, 143, 177, 175, 163, 131,  67,  63,  62,  74,  65,  36,  21, 115, 157, 152, 157, 154, 145, 147, 145, 139, 137, 141, 141, 138,
   177, 175, 178, 158,  65,  66,  61,  76, 143, 179, 175, 167, 169, 161, 171, 164, 160, 168, 182, 157, 176, 178, 164, 160, 164, 162, 171, 179, 168, 112,  48,  59,  58, 105, 108, 128,  69,  33,  89, 143, 152, 154, 149, 147, 147, 145, 138, 139, 143, 142,
   187, 183, 185, 166, 100, 100, 109, 115, 129, 166, 174, 165, 150, 160, 178, 148, 157, 164, 173, 164, 186, 183, 181, 165, 140, 131, 160, 181, 163,  99,  51,  60,  69, 112, 124, 152, 145,  69,  17,  65, 146, 153, 149, 141, 143, 143, 144, 142, 142, 139,
   186, 186, 186, 177, 116,  85,  83,  98, 130, 167, 154, 165, 167, 157, 148, 159, 162, 176, 179, 176, 181, 177, 170, 177, 169, 168, 169, 181, 147,  80,  66,  70, 107, 141, 136, 135, 150, 144,  46,  19,  82, 155, 149, 144, 147, 147, 145, 144, 143, 138,
   187, 186, 187, 179, 125, 113, 117, 114, 125, 171, 156, 148, 169, 156, 137, 160, 170, 180, 166, 181, 176, 169, 175, 180, 175, 173, 165, 185, 136,  41,  44,  89, 130, 133, 139, 152, 153, 156, 114,  26,  25,  97, 148, 147, 146, 147, 144, 142, 144, 143,
   188, 188, 190, 185, 145, 156, 137, 138, 176, 182, 173, 113, 121, 154, 151, 153, 162, 163, 164, 174, 167, 175, 168, 168, 133, 140, 143, 144, 103,  53,  25,  97, 148, 135, 144, 154, 150, 157, 154,  63,  22,  28, 115, 153, 142, 146, 142, 145, 142, 141,
   187, 186, 188, 192, 151, 155, 165, 164, 184, 185, 180, 153, 117, 154, 180, 161, 150, 155, 149, 155, 172, 174, 171, 152, 145, 103, 130, 132,  96,  63,  45,  92, 142, 129, 131, 143, 148, 162, 162, 124,  26,  21,  59, 148, 142, 146, 146, 148, 141, 138,
   191, 188, 185, 191, 163, 140, 168, 181, 179, 176, 177, 181, 151, 128, 162, 168, 154, 157, 154, 155, 169, 177, 176, 150, 157, 128, 134, 153, 128,  67,  80, 116, 138, 119, 115, 122, 136, 151, 158, 158,  57,  20,  30, 125, 145, 142, 142, 145, 143, 140,
   193, 191, 190, 192, 173, 134, 161, 178, 185, 193, 183, 180, 170, 130, 132, 181, 175, 158, 152, 158, 168, 177, 161, 139, 150, 126, 130, 135,  71,  91, 138, 141, 127, 144, 127, 117, 136, 142, 155, 155, 116,  23,  21,  87, 155, 146, 148, 147, 145, 142,
   192, 194, 197, 199, 183, 147, 157, 173, 184, 182, 184, 181, 173, 146, 106, 124, 165, 179, 156, 134, 156, 173, 161, 142, 147, 142, 118, 111,  79, 120, 153, 164, 137, 142, 124, 117, 124, 143, 148, 141, 154,  49,  20,  48, 146, 150, 148, 144, 142, 144,
   191, 191, 198, 198, 183, 154, 165, 172, 184, 188, 184, 174, 138, 155, 133, 110, 115, 154, 164, 157, 159, 167, 166, 172, 175, 160, 132,  93, 114, 140, 156, 178, 163, 134, 145, 115, 121, 138, 142, 140, 163,  99,  20,  25, 114, 147, 146, 141, 143, 141,
   192, 193, 197, 197, 188, 159, 165, 168, 182, 183, 195, 175, 154, 163, 156, 122, 114, 108, 134, 168, 160, 167, 170, 178, 185, 171, 149, 122, 120, 144, 164, 157, 149, 153, 148, 133, 126, 143, 141, 138, 156, 134,  29,  20,  98, 153, 146, 146, 148, 142,
   193, 194, 195, 194, 191, 165, 165, 169, 181, 192, 182, 164, 174, 187, 161, 135, 128, 106,  99, 132, 160, 182, 167, 164, 167, 170, 166, 132, 116, 147, 158, 146, 143, 133, 144, 138, 130, 129, 131, 144, 143, 146,  47,  14,  85, 156, 151, 150, 142, 145,
   194, 194, 197, 196, 190, 169, 156, 182, 185, 187, 187, 191, 180, 169, 163, 154, 149, 118, 117,  99, 142, 175, 166, 151, 164, 166, 160, 153, 136, 148, 124, 122, 151, 134, 138, 139, 130, 127, 140, 134, 128, 124,  94,  24,  82, 152, 150, 146, 144, 144,
   195, 195, 193, 194, 194, 170, 155, 181, 182, 181, 186, 186, 190, 158, 167, 160, 132, 123, 117,  94, 105, 149, 182, 152, 162, 167, 160, 159, 156, 120, 119, 122, 144, 137, 134, 138, 125, 132, 148, 138, 121, 116, 148,  86,  31, 137, 151, 147, 147, 143,
   195, 196, 192, 190, 191, 177, 151, 171, 181, 186, 189, 186, 166, 150, 172, 168, 146, 118, 128, 122, 116, 103, 153, 177, 164, 168, 160, 153, 147, 121, 119, 148, 166, 143, 128, 126, 140, 154, 144, 136, 121, 136, 148, 117,  20,  94, 157, 146, 148, 149,
   194, 194, 193, 191, 187, 173, 139, 161, 176, 180, 195, 181, 194, 180, 177, 170, 149, 138, 138, 139, 134, 130, 131, 169, 177, 178, 165, 156, 165, 144, 126, 125, 149, 155, 130, 136, 130, 137, 156, 129, 112, 143, 150, 139,  34,  45, 147, 147, 145, 146,
   194, 193, 189, 190, 192, 181,  86, 138, 169, 180, 186, 185, 176, 171, 203, 189, 141, 119, 111, 147, 130, 122, 143, 136, 160, 174, 170, 161, 169, 148, 156, 165, 147, 132, 129, 115, 134, 147, 149, 126, 115, 145, 151, 139,  42,  23, 126, 146, 145, 141,
   195, 191, 193, 191, 191, 197, 102,  91, 187, 175, 171, 183, 185, 175, 173, 164, 149, 141, 145, 154, 132, 147, 146, 151, 145, 154, 170, 155, 147, 152, 168, 157, 162, 144, 124, 106, 120, 141, 147, 125, 137, 141, 143, 149,  47,  16,  83, 146, 148, 147,
   194, 195, 193, 193, 192, 197, 142,  85, 183, 176, 176, 194, 180, 180, 184, 172, 160, 140, 175, 142, 131, 147, 146, 142, 150, 133, 145, 169, 145, 157, 156, 155, 151, 150, 122,  94, 122, 145, 154, 128, 133, 139, 148, 144,  48,  17,  51, 139, 145, 143,
   199, 196, 194, 194, 193, 194, 184, 135, 184, 183, 176, 193, 193, 183, 184, 172, 154, 159, 155, 121, 129, 141, 131, 110, 152, 158, 124, 146, 168, 164, 156, 161, 160, 132, 123,  85, 102, 144, 152, 130, 136, 150, 147, 136,  43,  17,  27, 120, 147, 147,
   196, 195, 196, 197, 196, 194, 198, 181, 178, 181, 182, 171, 184, 182, 176, 168, 161, 159, 164, 138, 144, 139, 130, 124, 131, 147, 147, 128, 145, 154, 149, 168, 169, 138, 122, 102,  85, 107, 140, 133, 145, 144, 140, 129,  36,  19,  18,  99, 147, 148,
   199, 199, 190, 194, 195, 195, 195, 193, 162, 176, 186, 150, 154, 164, 184, 173, 152, 155, 145, 134,  73,  83, 139, 132, 122, 143, 149, 155, 134, 146, 145, 159, 175, 137, 128, 134, 128,  41,  79, 118, 136, 143, 144, 114,  26,  21,  16,  85, 150, 144,
   200, 198, 194, 189, 191, 200, 193, 195, 180, 168, 178, 184, 159, 157, 167, 170, 175, 153, 126, 124,  88,  52,  95, 121, 129, 137, 153, 151, 149, 121, 131, 147, 164, 141, 127, 139, 146,  65,  52,  90, 118, 130, 130,  69,  16,  19,  17,  92, 152, 147,
   200, 197, 195, 195, 192, 196, 196, 192, 185, 151, 173, 196, 185, 189, 176, 153, 160, 147, 133, 132, 159,  86,  88, 116, 131, 133, 156, 164, 147, 143, 109, 134, 150, 142, 141, 147, 152,  43,  18,  73, 126, 110, 112,  30,  12,  16,  19, 113, 149, 150,
   196, 197, 197, 196, 191, 194, 193, 187, 189, 150, 169, 185, 188, 188, 154, 175, 168, 154, 152, 156, 152, 116,  93, 115, 128, 142, 169, 167, 164, 144, 124, 101, 114, 148, 140, 143, 161,  74,   8,  38, 116, 134, 116,  18,  13,  15,  25, 124, 146, 141,
   196, 195, 193, 193, 196, 192, 190, 187, 187, 180, 152, 174, 182, 172, 170, 168, 169, 171, 181, 194, 169, 174, 150, 133, 133, 132, 161, 164, 168, 155, 151, 133,  82,  91, 134, 128, 148, 123,  14,  40, 130, 152, 107,  21,  14,  14,  50, 142, 141, 144,
   198, 195, 195, 195, 195, 193, 190, 189, 186, 192, 161, 174, 181, 176, 178, 182, 174, 172, 177, 177, 176, 176, 173, 167, 163, 143, 162, 157, 154, 147, 159, 166, 129,  80,  81, 129, 128, 148,  89,  47,  98, 133,  71,  21,  16,  17,  97, 149, 142, 148,
   197, 200, 196, 197, 191, 193, 190, 189, 190, 188, 178, 159, 184, 186, 176, 169, 174, 179, 183, 153, 176, 153, 168, 183, 169, 158, 153, 151, 145, 144, 149, 157, 157, 122,  71,  65, 119, 129, 139, 101, 109, 126,  33,  22,  17,  30, 132, 145, 145, 145,
   193, 195, 196, 193, 192, 193, 190, 190, 186, 188, 189, 160, 157, 179, 178, 167, 175, 183, 169, 172, 167, 159, 173, 174, 173, 165, 151, 150, 149, 144, 151, 153, 151, 159, 119,  63,  56, 104, 115, 118, 117, 126,  58,  22,  16,  55, 144, 147, 150, 142,
   194, 196, 197, 193, 194, 191, 191, 189, 185, 189, 189, 184, 156, 176, 189, 168, 173, 176, 170, 178, 167, 158, 153, 150, 168, 163, 164, 148, 138, 142, 158, 165, 160, 155, 162, 129,  78,  54,  77,  80, 109, 112,  90,  22,  16, 101, 149, 147, 147, 141,
   192, 197, 193, 191, 191, 191, 189, 192, 187, 188, 191, 189, 176, 145, 168, 179, 179, 183, 173, 175, 161, 157, 153, 157, 172, 170, 157, 157, 149, 140, 140, 144, 153, 158, 148, 144, 131,  91,  56,  50,  64,  77,  88,  62, 108, 143, 145, 144, 145, 143,
   193, 195, 192, 190, 192, 191, 192, 188, 187, 186, 186, 190, 184, 165, 145, 169, 172, 169, 160, 157, 144, 141, 158, 151, 159, 153, 143, 148, 138, 134, 148, 125, 153, 165, 159, 157, 156, 139, 110,  73,  45,  29,  16,  31, 119, 151, 147, 147, 144, 147,
   193, 192, 191, 193, 193, 190, 190, 190, 187, 181, 184, 182, 189, 187, 170, 166, 172, 155, 162, 158, 154, 153, 153, 159, 155, 147, 151, 167, 137, 134, 146, 130, 152, 161, 167, 155, 140, 140, 141, 109,  67,  40,  26,   8,  24,  98, 143, 149, 146, 144,
   194, 191, 193, 194, 192, 194, 192, 193, 189, 186, 191, 184, 178, 183, 187, 180, 177, 169, 175, 163, 178, 165, 155, 152, 151, 150, 144, 157, 128, 144, 126, 129, 147, 151, 143, 133, 114, 128, 133, 137, 112,  65,  43,  25,  12,  17,  97, 151, 154, 153,
   195, 195, 194, 194, 198, 194, 188, 189, 187, 190, 187, 187, 184, 184, 194, 194, 188, 182, 169, 170, 145, 175, 160, 144, 141, 152, 152, 137, 140, 146, 124, 159, 142, 132, 129, 126, 129, 137, 131, 133, 141,  96,  59,  51,  19,  14, 104, 152, 101,  91,
   193, 191, 190, 192, 196, 195, 189, 185, 193, 194, 188, 191, 189, 189, 189, 186, 182, 185, 179, 178, 160, 177, 160, 143, 142, 151, 141, 140, 145, 136, 142, 153, 136, 137, 150, 134, 136, 140, 130, 119, 118,  55,  38,  97,  76,  33, 132, 159,  81,  15,
   193, 190, 195, 196, 189, 190, 188, 185, 189, 188, 185, 179, 184, 193, 187, 178, 182, 181, 184, 181, 182, 176, 168, 157, 154, 151, 151, 143, 134, 143, 135, 127, 120, 126, 145, 146, 139, 128, 114,  99,  82,  64,  85, 156, 155,  91, 136, 156,  76,  37,
   194, 194, 193, 194, 192, 196, 198, 192, 190, 189, 187, 185, 191, 189, 188, 190, 187, 183, 185, 180, 177, 189, 186, 172, 177, 173, 159, 142, 143, 139, 120, 124, 127, 149, 161, 159, 157, 157, 153, 151, 153, 160, 161, 159, 174, 116, 105, 150, 113, 126,
   192, 195, 195, 193, 190, 193, 189, 190, 193, 192, 192, 189, 190, 186, 183, 183, 183, 181, 184, 180, 177, 185, 186, 182, 182, 180, 181, 175, 173, 167, 167, 166, 171, 164, 165, 165, 161, 165, 162, 161, 161, 160, 151, 150, 161, 149, 124, 148, 152, 144,
   194, 192, 194, 194, 192, 191, 189, 190, 192, 187, 187, 194, 189, 181, 178, 176, 182, 181, 187, 185, 181, 183, 185, 181, 185, 185, 180, 182, 177, 173, 172, 172, 168, 169, 167, 164, 163, 167, 164, 166, 165, 154, 151, 151, 149, 151, 148, 147, 145, 138,
   197, 193, 192, 188, 191, 195, 192, 189, 182, 188, 189, 188, 193, 181, 183, 175, 178, 184, 187, 187, 183, 187, 182, 181, 177, 180, 178, 173, 173, 171, 175, 171, 167, 168, 172, 173, 166, 161, 162, 162, 163, 160, 151, 151, 151, 151, 147, 143, 140, 136
};

B = '{
 184, 180, 186, 182, 180, 177, 178, 179, 177, 177, 171, 173, 173, 170, 173, 174, 171, 172, 171, 164, 165, 167, 169, 161, 162, 162, 167, 157, 151, 153, 162, 166, 166, 152, 146, 154, 152, 163, 156, 145, 154, 151, 147, 152, 146, 141, 135, 134, 141, 136,
   187, 188, 187, 180, 182, 178, 177, 177, 175, 177, 176, 174, 171, 168, 173, 171, 168, 170, 171, 162, 166, 164, 169, 155, 163, 161, 160, 153, 157, 156, 155, 160, 162, 158, 154, 157, 155, 159, 156, 149, 148, 148, 145, 147, 147, 144, 138, 139, 139, 143,
   188, 189, 185, 180, 180, 179, 176, 178, 179, 178, 181, 177, 172, 174, 176, 168, 165, 174, 170, 163, 168, 168, 167, 159, 164, 167, 166, 165, 155, 159, 157, 160, 156, 157, 158, 154, 158, 156, 161, 154, 153, 151, 150, 146, 145, 152, 144, 142, 137, 136,
   190, 184, 179, 179, 184, 189, 184, 180, 179, 179, 178, 170, 164, 165, 165, 164, 160, 160, 164, 158, 163, 158, 153, 159, 158, 172, 159, 160, 162, 157, 156, 157, 156, 154, 152, 157, 154, 151, 150, 154, 155, 150, 150, 147, 144, 147, 147, 143, 141, 134,
   189, 184, 185, 187, 148, 146, 171, 179, 166, 153, 135, 108,  91,  86,  83,  95,  88,  80,  95, 104, 113, 113, 108,  97,  75,  68,  79, 103,  99, 110, 134, 154, 159, 155, 155, 161, 162, 156, 146, 151, 156, 156, 148, 145, 144, 145, 144, 143, 142, 140,
   184, 184, 186, 158,  54,  19,  33,  59,  30,  50,  95, 101, 115, 105,  90,  97,  95,  96,  96, 118, 108,  98, 111, 101,  96,  92,  63,  34,  27,  35,  41,  50,  62,  96, 142, 160, 158, 151, 152, 148, 150, 159, 154, 148, 147, 142, 145, 148, 142, 143,
   187, 185, 184,  89,  24,  12,   9,  23,  46,  56, 124, 131, 128, 130, 122, 129, 134, 133, 125, 137, 121, 113, 132, 130, 108,  93,  93,  96,  65,  28,  29,  29,  30,  28,  49, 108, 150, 159, 155, 150, 157, 156, 155, 151, 144, 145, 144, 142, 146, 144,
   189, 190, 184,  67,  10,  18,  41,  64, 105, 117, 113, 134, 125, 130, 144, 131, 129, 120, 135, 139, 106, 104, 138, 144, 124, 101, 100,  97,  98,  74,  30,  16,  21,  25,  25,  28,  68, 151, 161, 157, 164, 163, 155, 149, 144, 146, 143, 144, 146, 143,
   188, 182, 186, 129,  13,  26,  26,  65, 101, 127, 115, 131, 108, 116, 139, 140, 124, 138, 150, 131, 123, 124, 110, 128, 140, 120, 123, 111, 100,  73,  13,  12,  13,  25,  27,  26,  28, 121, 163, 158, 162, 158, 152, 155, 151, 145, 143, 147, 147, 144,
   184, 181, 185, 142,  15,  20,  24,  45, 100, 123, 122, 123, 127, 108, 126, 130, 125, 122, 144, 121, 145, 147, 127, 105, 131, 138, 121, 126, 115,  67,   5,  16,  15,  46,  44,  73,  41,  26,  88, 147, 153, 157, 155, 154, 153, 151, 144, 147, 150, 149,
   193, 189, 193, 143,  14,  23,  32,  62,  97, 127, 127, 121, 111, 108, 138, 125, 134, 118, 130, 125, 146, 144, 144, 112, 104, 112, 113, 122,  99,  37,   8,  16,  19,  53,  60,  93,  93,  35,   9,  66, 146, 154, 154, 148, 149, 149, 150, 150, 151, 147,
   192, 192, 195, 166,  42,  31,  41,  70, 105, 136, 108, 117, 130, 110, 115, 130, 128, 132, 137, 136, 142, 137, 136, 135, 119, 134, 119, 115,  81,  30,  21,  23,  52,  85,  81,  76,  88,  93,  21,  11,  80, 157, 154, 151, 153, 153, 152, 152, 151, 146,
   192, 191, 194, 174,  58,  57,  89,  94, 100, 140, 115, 105, 132, 116, 101, 116, 124, 140, 126, 145, 143, 132, 142, 141, 129, 124, 115, 133,  89,  24,  18,  43,  79,  87,  98,  94,  93, 104,  63,   7,  16,  94, 151, 153, 151, 152, 149, 149, 151, 150,
   192, 192, 196, 186,  88,  91, 102, 105, 136, 142, 137,  80,  85, 117, 110, 106, 118, 126, 121, 136, 134, 135, 129, 131, 111, 110, 111, 119,  80,  45,  19,  66, 100,  83,  99, 103,  94, 105,  94,  33,   8,  20, 114, 158, 146, 150, 147, 151, 147, 147,
   191, 190, 193, 195, 101,  89, 116, 121, 141, 140, 138, 117,  77, 110, 139, 118, 103, 111, 108, 113, 140, 137, 130, 124, 135,  90, 113, 120,  83,  52,  31,  60,  92,  80,  88,  93,  97, 114, 113,  76,   5,  10,  55, 149, 146, 149, 150, 154, 147, 145,
   195, 192, 190, 198, 123,  73, 118, 141, 144, 138, 141, 150, 112,  75, 116, 132, 111, 111, 109, 111, 138, 144, 139, 127, 144, 112, 118, 142, 114,  46,  54,  71,  82,  94,  73,  68,  86, 106, 111,  96,  25,   8,  20, 125, 148, 146, 147, 150, 148, 146,
   197, 195, 194, 200, 144,  65, 108, 136, 150, 161, 155, 151, 134,  76,  80, 147, 140, 121, 106, 118, 138, 142, 123, 123, 139, 114, 116, 123,  61,  63,  99,  94,  66, 110,  71,  64,  89,  99, 105,  92,  64,   5,   6,  86, 157, 151, 156, 151, 148, 146,
   196, 198, 200, 206, 161,  82, 104, 128, 141, 141, 145, 140, 138, 102,  53,  76, 123, 146, 120,  98, 125, 137, 128, 123, 131, 127,  93,  93,  60,  78, 100, 118,  80,  87,  69,  65,  73,  97, 101,  84,  93,  18,   3,  44, 148, 154, 155, 149, 146, 148,
   195, 195, 201, 205, 167,  93, 108, 122, 137, 146, 148, 142, 115, 122,  84,  55,  66, 115, 127, 124, 127, 129, 129, 143, 145, 126,  92,  64,  72,  87, 109, 137, 116,  80,  92,  57,  61,  85,  94,  88, 103,  54,   3,  16, 115, 150, 151, 145, 147, 145,
   196, 197, 200, 202, 178, 106, 105, 115, 139, 147, 165, 159, 138, 133, 114,  77,  69,  59,  86, 132, 126, 132, 132, 149, 151, 123, 100,  70,  68,  95, 112,  98,  97,  99,  99,  81,  75,  90,  87,  85, 103,  79,   6,  10,  94, 153, 148, 150, 152, 146,
   197, 198, 198, 199, 188, 115, 109, 121, 137, 157, 155, 142, 144, 148, 122,  93,  81,  51,  43,  86, 121, 146, 126, 130, 130, 126, 121,  84,  71,  97, 110, 100,  95,  73,  95,  90,  83,  77,  74,  87,  84,  89,  15,   7,  81, 156, 152, 154, 146, 149,
   198, 198, 200, 202, 194, 123, 105, 139, 144, 151, 149, 148, 142, 139, 130, 117, 109,  72,  63,  38,  91, 134, 124, 115, 123, 126, 119, 109,  84,  95,  93, 103, 117,  81,  87,  86,  76,  72,  85,  77,  76,  84,  46,   9,  78, 152, 152, 150, 148, 148,
   199, 199, 197, 197, 201, 136,  98, 138, 147, 150, 140, 137, 153, 127, 138, 125,  90,  76,  67,  42,  47,  98, 144, 118, 123, 131, 118, 116, 110,  78,  98, 103,  97,  94,  89,  89,  71,  79,  99,  88,  72,  80,  90,  46,  21, 135, 157, 151, 151, 147,
   199, 200, 196, 193, 198, 157,  89, 116, 141, 150, 147, 145, 127, 113, 144, 139, 111,  71,  76,  74,  57,  38, 104, 139, 132, 128, 110, 105, 118,  99, 101, 115, 114,  98,  78,  79,  96, 106,  90,  80,  62,  81,  85,  69,   1,  91, 159, 150, 152, 153,
   198, 198, 197, 193, 194, 165,  83, 105, 137, 141, 157, 147, 158, 145, 145, 142, 125, 110, 104,  98,  88,  73,  74, 113, 130, 139, 118, 113, 145, 132, 102,  83,  99, 106,  70,  86,  96, 101, 110,  82,  58,  86,  93,  87,   7,  42, 146, 151, 149, 151,
   198, 197, 194, 195, 195, 180,  67, 102, 127, 138, 149, 151, 135, 131, 178, 180, 132, 107,  89, 111,  86,  75,  92,  70, 100, 129, 128, 122, 149, 133, 116, 115,  99,  73,  64,  59,  92, 106, 102,  78,  62,  93,  98,  78,  11,  16, 122, 148, 149, 148,
   199, 195, 197, 197, 194, 197,  99,  72, 153, 136, 133, 147, 150, 138, 147, 154, 139, 128, 123, 122,  95, 111, 107, 103,  95,  93, 113, 116, 128, 130, 127, 110, 117,  92,  67,  52,  74,  93,  94,  69,  80,  89,  89,  87,  16,   8,  78, 147, 153, 155,
   198, 199, 197, 198, 195, 197, 141,  68, 146, 136, 134, 156, 153, 149, 152, 147, 134, 116, 146, 106,  94, 109, 100,  97,  98,  61,  67, 114, 110, 114, 107, 102, 100,  96,  68,  43,  72,  95, 105,  77,  78,  87,  95,  82,  16,   8,  45, 141, 149, 150,
   201, 199, 196, 198, 197, 198, 184,  96, 143, 141, 130, 155, 165, 152, 153, 140, 125, 142, 135,  91,  81,  84,  91,  79, 112, 105,  60,  80, 108, 107, 103, 107, 107,  73,  62,  29,  49,  93,  99,  75,  83, 100,  92,  73,  12,   9,  21, 121, 148, 149,
   198, 197, 198, 201, 200, 198, 198, 144, 127, 135, 142, 139, 153, 145, 141, 135, 136, 145, 148, 117, 114, 103, 105, 108, 106, 101,  91,  65,  75,  91,  96, 122, 123,  86,  65,  45,  38,  66,  84,  75,  91,  92,  83,  68,  10,   9,  12, 100, 148, 149,
   201, 201, 192, 198, 199, 199, 200, 177, 107, 131, 154, 127, 123, 125, 142, 137, 131, 143, 130, 119,  61,  69, 118, 116,  99,  96,  94,  97,  70,  83,  87, 110, 130,  86,  76,  75,  84,  25,  45,  64,  80,  87,  85,  57,   6,   8,  11,  86, 151, 145,
   202, 200, 196, 191, 193, 202, 196, 192, 133, 118, 139, 156, 131, 120, 124, 139, 159, 143, 110, 107,  75,  40,  74,  95, 105,  95,  98,  99,  99,  66,  73,  89, 108,  85,  75,  83, 105,  47,  29,  50,  56,  77,  71,  30,   3,   9,  12,  92, 154, 150,
   202, 199, 197, 197, 194, 197, 195, 203, 151,  97, 138, 166, 148, 154, 139, 113, 134, 131, 117, 112, 142,  73,  72,  99, 116, 103, 105, 111, 100,  88,  44,  69,  86,  79,  84,  94, 111,  25,   8,  50,  73,  69,  58,   8,   5,  11,  16, 112, 152, 154,
   198, 199, 199, 198, 193, 197, 196, 193, 180,  96, 127, 154, 156, 148, 112, 144, 136, 116, 121, 133, 127,  88,  65,  96, 108, 103, 112, 111, 108,  85,  61,  35,  49,  81,  80,  92, 117,  48,   3,  27,  74,  86,  53,   2,   8,  12,  23, 124, 148, 145,
   198, 197, 195, 195, 198, 194, 194, 187, 193, 143,  90, 136, 144, 125, 129, 144, 135, 127, 143, 167, 132, 134,  95,  79,  79,  76, 108, 115, 121, 111, 110,  77,  18,  32,  77,  69,  98,  88,   2,  25,  79,  90,  34,   5,   8,  10,  52, 143, 143, 146,
   200, 197, 197, 197, 197, 195, 193, 193, 192, 184, 104, 125, 146, 135, 143, 147, 135, 138, 147, 143, 137, 138, 131, 124, 115,  90, 118, 111, 107, 102, 115, 121,  76,  21,  23,  71,  69,  98,  53,  18,  60,  77,  20,   7,   7,  11, 100, 151, 144, 150,
   199, 202, 198, 199, 193, 195, 194, 194, 195, 191, 145,  97, 148, 155, 143, 130, 136, 148, 150, 110, 139, 113, 130, 151, 124, 111, 111, 104,  95,  95, 100, 113, 117,  73,  19,  18,  63,  69,  84,  54,  65,  76,  15,   8,   7,  25, 135, 147, 147, 147,
   195, 197, 198, 196, 195, 197, 194, 193, 189, 190, 183, 112, 104, 139, 143, 130, 146, 155, 129, 131, 131, 115, 128, 133, 132, 126, 110, 102,  99,  98, 107, 109, 112, 120,  70,  12,   9,  50,  67,  72,  61,  76,  38,   8,   5,  49, 145, 148, 152, 145,
   196, 198, 199, 197, 198, 195, 193, 191, 187, 193, 195, 173, 128, 145, 155, 133, 127, 130, 135, 153, 134, 111, 109, 109, 135, 127, 125, 109,  94,  96, 110, 118, 113, 108, 108,  74,  26,   4,  30,  38,  59,  56,  51,   4,   8,  96, 148, 147, 150, 146,
   194, 199, 195, 194, 195, 195, 191, 194, 189, 190, 195, 195, 174, 110, 115, 142, 143, 146, 145, 144, 127, 112, 115, 123, 135, 133, 119, 118, 102,  89,  86,  91, 101, 106, 101,  98,  82,  44,  11,  11,  27,  32,  55,  46, 106, 143, 145, 144, 147, 147,
   195, 197, 194, 193, 196, 195, 194, 191, 190, 190, 189, 194, 187, 135,  92, 132, 143, 139, 113, 111,  99,  92, 111, 111, 113, 106,  97, 102,  92,  87, 104,  83, 108, 121, 121, 120, 113,  93,  63,  27,   9,   9,   5,  29, 121, 154, 148, 148, 146, 150,
   195, 194, 193, 197, 197, 194, 194, 194, 191, 185, 188, 186, 193, 183, 143, 123, 131, 117, 123, 122, 112, 105, 107, 119, 111,  99, 108, 129,  99,  94, 104,  89, 110, 128, 133, 119, 100,  94, 101,  67,  19,   7,  13,   6,  27, 104, 146, 150, 147, 146,
   196, 193, 195, 198, 196, 198, 196, 197, 193, 190, 195, 188, 180, 190, 190, 157, 136, 128, 140, 133, 142, 125, 120, 120, 111, 113, 106, 118,  82, 104,  81,  80, 106, 117, 101,  88,  70,  85,  96,  98,  59,  13,  12,   8,   8,  20, 102, 151, 153, 151,
   197, 197, 196, 197, 201, 197, 191, 192, 190, 194, 191, 191, 190, 185, 196, 202, 182, 159, 136, 129, 101, 130, 128, 107,  97, 111, 112,  95,  90, 103,  76, 110,  99,  87,  80,  76,  83,  96,  94,  93,  87,  45,  20,  10,   3,  17,  97, 134,  88,  88,
   195, 193, 192, 194, 198, 197, 191, 187, 195, 197, 192, 195, 193, 193, 193, 193, 192, 187, 175, 169, 134, 130, 111,  92, 100, 108,  98,  98, 102,  86,  96, 101,  74,  79,  99,  82,  92, 103,  90,  77,  70,  26,  20,  43,  25,  20,  89,  91,  38,  10,
   195, 192, 197, 198, 191, 192, 190, 187, 191, 191, 189, 183, 188, 197, 190, 183, 188, 184, 186, 188, 183, 162, 138, 111, 103,  95, 100,  97,  84,  88,  84,  71,  64,  75,  88,  82,  82,  82,  75,  68,  62,  61,  81, 123,  77,  24,  71,  81,  37,  32,
   197, 197, 195, 196, 194, 198, 201, 195, 192, 192, 191, 190, 195, 193, 192, 193, 189, 187, 190, 187, 187, 193, 189, 166, 168, 150, 124,  98,  94,  86,  72,  85, 106, 138, 143, 129, 122, 130, 138, 147, 153, 160, 162, 155, 124,  43,  61, 109,  98, 129,
   195, 199, 199, 195, 192, 195, 192, 194, 196, 196, 196, 193, 195, 192, 189, 188, 187, 184, 189, 187, 183, 190, 190, 187, 188, 184, 184, 177, 171, 164, 164, 166, 173, 167, 168, 168, 163, 166, 164, 164, 163, 160, 153, 152, 151, 128, 120, 147, 152, 144,
   198, 196, 198, 196, 194, 193, 193, 194, 196, 192, 191, 198, 194, 187, 185, 182, 186, 185, 192, 191, 187, 188, 189, 185, 189, 189, 184, 187, 180, 176, 175, 175, 170, 171, 169, 167, 165, 169, 166, 168, 166, 155, 152, 151, 153, 160, 149, 149, 147, 140,
   201, 197, 196, 190, 193, 196, 195, 193, 186, 192, 193, 192, 198, 187, 189, 180, 182, 188, 192, 194, 189, 193, 186, 185, 181, 184, 182, 177, 177, 175, 179, 175, 171, 172, 175, 175, 168, 163, 164, 164, 165, 161, 152, 155, 158, 153, 155, 148, 144, 140
};
wr_en = 0;
reset = 1;
#20;
reset = 0;
#20;
@(posedge clk_100);
//150 * 150 = 2500 for features verifiation
for(i = 0;i<2500;i++)
begin
    b <= B[i];
    g <= G[i];
    r <= R[i];
    wr_en <= 1;
    @(posedge clk_100);
    wr_en <= 0;
    @(posedge clk_100);
    repeat(100) begin
        @(posedge clk_100);
    end
end

end


always begin
#4 clk_100 = ~clk_100;
end

    
endmodule
