`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/14/2022 11:32:31 PM
// Design Name: 
// Module Name: Fix_NN
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/11/2022 12:03:41 AM
// Design Name: 
// Module Name: Fix_NN
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Fix_NN(
input clk,reset,start_fix_conv,
input [31:0]LBP_161, LBP_156, LBP_137, LBP_136, LBP_132, LBP_128, LBP_125, LBP_43, LBP_38, 
LBP_32, LBP_25, LBP_19, LBP_14, LBP_7,
input [31:0]a_bin198 , a_bin199, b_bin208,
output reg [2:0]EB_LB_HD = 0,
output reg NN_done = 0
);

reg [7:0]EB_count=0,HD_count=0,LB_count=0;

reg [29:0] w8_L1_N1_0= 30'h00000000,  w8_L1_N1_1= 30'h00000000,  w8_L1_N1_2= 30'h00000000,  w8_L1_N1_3= 30'h00000000,  w8_L1_N1_4= 30'h00000000,  w8_L1_N1_5= 30'h00000000,  w8_L1_N1_6= 30'h00000000,  w8_L1_N1_7= 30'h00000000,  w8_L1_N1_8= 30'h00000000,  w8_L1_N1_9= 30'h00000000,  w8_L1_N1_10= 30'h00000000,  w8_L1_N1_11= 30'h00000000,  w8_L1_N1_12= 30'h00000000,  w8_L1_N1_13= 30'h00000000,  w8_L1_N1_14= 30'h00000000,  w8_L1_N1_15= 30'h00000000,  w8_L1_N1_16= 30'h00000000;
reg [29:0] w8_L1_N2_0= 30'h00000000,  w8_L1_N2_1= 30'h00000000,  w8_L1_N2_2= 30'h00000000,  w8_L1_N2_3= 30'h00000000,  w8_L1_N2_4= 30'h00000000,  w8_L1_N2_5= 30'h00000000,  w8_L1_N2_6= 30'h00000000,  w8_L1_N2_7= 30'h00000000,  w8_L1_N2_8= 30'h00000000,  w8_L1_N2_9= 30'h00000000,  w8_L1_N2_10= 30'h00000000,  w8_L1_N2_11= 30'h00000000,  w8_L1_N2_12= 30'h00000000,  w8_L1_N2_13= 30'h00000000,  w8_L1_N2_14= 30'h00000000,  w8_L1_N2_15= 30'h00000000,  w8_L1_N2_16= 30'h00000000;
reg [29:0] w8_L1_N3_0= 30'h3ffff0d2,  w8_L1_N3_1= 30'h3fff7ac9,  w8_L1_N3_2= 30'h0002b936,  w8_L1_N3_3= 30'h3ff89575,  w8_L1_N3_4= 30'h3ff5a418,  w8_L1_N3_5= 30'h3ffa217d,  w8_L1_N3_6= 30'h3ff64666,  w8_L1_N3_7= 30'h3ff65c18,  w8_L1_N3_8= 30'h3ff6aaf1,  w8_L1_N3_9= 30'h3ff5801c,  w8_L1_N3_10= 30'h3ff8abc6,  w8_L1_N3_11= 30'h3ff583ad,  w8_L1_N3_12= 30'h3ff95d85,  w8_L1_N3_13= 30'h3ff642fb,  w8_L1_N3_14= 30'h3ffa0229,  w8_L1_N3_15= 30'h3ff60879,  w8_L1_N3_16= 30'h3ff4f587;
reg [29:0] w8_L1_N4_0= 30'h0002cad5,  w8_L1_N4_1= 30'h3ffeb8ee,  w8_L1_N4_2= 30'h0002c08b,  w8_L1_N4_3= 30'h3febb6f4,  w8_L1_N4_4= 30'h3fe90f01,  w8_L1_N4_5= 30'h3fee7a7e,  w8_L1_N4_6= 30'h3fe61acb,  w8_L1_N4_7= 30'h3fecb101,  w8_L1_N4_8= 30'h3fe86c86,  w8_L1_N4_9= 30'h3fea2747,  w8_L1_N4_10= 30'h3fecd3c0,  w8_L1_N4_11= 30'h3fea4d27,  w8_L1_N4_12= 30'h3fedf4d0,  w8_L1_N4_13= 30'h3feb4ea5,  w8_L1_N4_14= 30'h3fef4763,  w8_L1_N4_15= 30'h3fe9d57f,  w8_L1_N4_16= 30'h3feae944;
reg [29:0] w8_L1_N5_0= 30'h00000000,  w8_L1_N5_1= 30'h00000000,  w8_L1_N5_2= 30'h000002ca,  w8_L1_N5_3= 30'h00000000,  w8_L1_N5_4= 30'h00000000,  w8_L1_N5_5= 30'h00000000,  w8_L1_N5_6= 30'h00000000,  w8_L1_N5_7= 30'h00000000,  w8_L1_N5_8= 30'h00000000,  w8_L1_N5_9= 30'h00000000,  w8_L1_N5_10= 30'h00000000,  w8_L1_N5_11= 30'h00000000,  w8_L1_N5_12= 30'h00000000,  w8_L1_N5_13= 30'h00000000,  w8_L1_N5_14= 30'h00000000,  w8_L1_N5_15= 30'h00000000,  w8_L1_N5_16= 30'h00000000;
reg [29:0] w8_L1_N6_0= 30'h00000000,  w8_L1_N6_1= 30'h00000000,  w8_L1_N6_2= 30'h00000000,  w8_L1_N6_3= 30'h00000000,  w8_L1_N6_4= 30'h00000000,  w8_L1_N6_5= 30'h00000000,  w8_L1_N6_6= 30'h00000000,  w8_L1_N6_7= 30'h00000000,  w8_L1_N6_8= 30'h00000000,  w8_L1_N6_9= 30'h00000000,  w8_L1_N6_10= 30'h00000000,  w8_L1_N6_11= 30'h00000000,  w8_L1_N6_12= 30'h00000000,  w8_L1_N6_13= 30'h00000000,  w8_L1_N6_14= 30'h00000000,  w8_L1_N6_15= 30'h00000000,  w8_L1_N6_16= 30'h00000000;
reg [29:0] w8_L1_N7_0= 30'h00000000,  w8_L1_N7_1= 30'h00000000,  w8_L1_N7_2= 30'h00000000,  w8_L1_N7_3= 30'h00000000,  w8_L1_N7_4= 30'h00000000,  w8_L1_N7_5= 30'h00000000,  w8_L1_N7_6= 30'h00000000,  w8_L1_N7_7= 30'h00000000,  w8_L1_N7_8= 30'h00000000,  w8_L1_N7_9= 30'h00000000,  w8_L1_N7_10= 30'h00000000,  w8_L1_N7_11= 30'h00000000,  w8_L1_N7_12= 30'h00000000,  w8_L1_N7_13= 30'h00000000,  w8_L1_N7_14= 30'h00000000,  w8_L1_N7_15= 30'h00000000,  w8_L1_N7_16= 30'h00000000;
reg [29:0] w8_L1_N8_0= 30'h3ffbbe40,  w8_L1_N8_1= 30'h00015c80,  w8_L1_N8_2= 30'h3ffe5bdb,  w8_L1_N8_3= 30'h00173835,  w8_L1_N8_4= 30'h001af78c,  w8_L1_N8_5= 30'h00155c5a,  w8_L1_N8_6= 30'h001e8afb,  w8_L1_N8_7= 30'h00187cc9,  w8_L1_N8_8= 30'h001be793,  w8_L1_N8_9= 30'h00186d22,  w8_L1_N8_10= 30'h0016cd7d,  w8_L1_N8_11= 30'h00198ebb,  w8_L1_N8_12= 30'h00162149,  w8_L1_N8_13= 30'h00174fec,  w8_L1_N8_14= 30'h0016466b,  w8_L1_N8_15= 30'h0019efee,  w8_L1_N8_16= 30'h00184e40;
reg [29:0] w8_L1_N9_0= 30'h0004ffd5,  w8_L1_N9_1= 30'h00044ecf,  w8_L1_N9_2= 30'h3ffdccdb,  w8_L1_N9_3= 30'h3fe87742,  w8_L1_N9_4= 30'h3fe6848a,  w8_L1_N9_5= 30'h3fe9549e,  w8_L1_N9_6= 30'h3fdfd93e,  w8_L1_N9_7= 30'h3fe7bbd6,  w8_L1_N9_8= 30'h3fe333c1,  w8_L1_N9_9= 30'h3fe4f65b,  w8_L1_N9_10= 30'h3fe88c9b,  w8_L1_N9_11= 30'h3fe6c235,  w8_L1_N9_12= 30'h3fe9a6b3,  w8_L1_N9_13= 30'h3fe77f5f,  w8_L1_N9_14= 30'h3fe9db52,  w8_L1_N9_15= 30'h3fe5da8d,  w8_L1_N9_16= 30'h3fe63688;
reg [29:0] w8_L1_N10_0= 30'h3ffe2669,  w8_L1_N10_1= 30'h00015932,  w8_L1_N10_2= 30'h000083bc,  w8_L1_N10_3= 30'h000e4326,  w8_L1_N10_4= 30'h0011f1bf,  w8_L1_N10_5= 30'h000cd998,  w8_L1_N10_6= 30'h0012aec6,  w8_L1_N10_7= 30'h00103e6b,  w8_L1_N10_8= 30'h0011ff75,  w8_L1_N10_9= 30'h0011cd64,  w8_L1_N10_10= 30'h000f35f9,  w8_L1_N10_11= 30'h00122a67,  w8_L1_N10_12= 30'h000de61d,  w8_L1_N10_13= 30'h000f76c0,  w8_L1_N10_14= 30'h000c888f,  w8_L1_N10_15= 30'h0010d337,  w8_L1_N10_16= 30'h00110363;
reg [29:0] w8_L1_N11_0= 30'h3ffe416b,  w8_L1_N11_1= 30'h0000d39e,  w8_L1_N11_2= 30'h3ffd526f,  w8_L1_N11_3= 30'h00161024,  w8_L1_N11_4= 30'h001b3ae9,  w8_L1_N11_5= 30'h0014fd13,  w8_L1_N11_6= 30'h001c8a33,  w8_L1_N11_7= 30'h001a0af2,  w8_L1_N11_8= 30'h001b43e6,  w8_L1_N11_9= 30'h001a7646,  w8_L1_N11_10= 30'h001677d3,  w8_L1_N11_11= 30'h001acf98,  w8_L1_N11_12= 30'h001695e0,  w8_L1_N11_13= 30'h0019308c,  w8_L1_N11_14= 30'h00153da8,  w8_L1_N11_15= 30'h001953d7,  w8_L1_N11_16= 30'h0019f7f9;
reg [29:0] w8_L1_N12_0= 30'h00000000,  w8_L1_N12_1= 30'h00000000,  w8_L1_N12_2= 30'h00000000,  w8_L1_N12_3= 30'h00000000,  w8_L1_N12_4= 30'h00000000,  w8_L1_N12_5= 30'h00000000,  w8_L1_N12_6= 30'h00000000,  w8_L1_N12_7= 30'h00000000,  w8_L1_N12_8= 30'h00000000,  w8_L1_N12_9= 30'h00000000,  w8_L1_N12_10= 30'h00000000,  w8_L1_N12_11= 30'h00000000,  w8_L1_N12_12= 30'h00000000,  w8_L1_N12_13= 30'h00000000,  w8_L1_N12_14= 30'h00000000,  w8_L1_N12_15= 30'h00000000,  w8_L1_N12_16= 30'h00000000;
reg [29:0] w8_L1_N13_0= 30'h3fffbdf7,  w8_L1_N13_1= 30'h0000415f,  w8_L1_N13_2= 30'h0003a7e8,  w8_L1_N13_3= 30'h3ff89c8e,  w8_L1_N13_4= 30'h3ff656a9,  w8_L1_N13_5= 30'h3ffa3cc3,  w8_L1_N13_6= 30'h3ff6b206,  w8_L1_N13_7= 30'h3ff65ace,  w8_L1_N13_8= 30'h3ff73ca3,  w8_L1_N13_9= 30'h3ff56438,  w8_L1_N13_10= 30'h3ff8b319,  w8_L1_N13_11= 30'h3ff61b73,  w8_L1_N13_12= 30'h3ff94d71,  w8_L1_N13_13= 30'h3ff741e8,  w8_L1_N13_14= 30'h3ffa5e9b,  w8_L1_N13_15= 30'h3ff6b2f6,  w8_L1_N13_16= 30'h3ff5d027;
reg [29:0] w8_L1_N14_0= 30'h3ffedf64,  w8_L1_N14_1= 30'h000577d8,  w8_L1_N14_2= 30'h3fff2f97,  w8_L1_N14_3= 30'h3ffb3536,  w8_L1_N14_4= 30'h3ffad52a,  w8_L1_N14_5= 30'h3ffbf9c0,  w8_L1_N14_6= 30'h3ff73bc4,  w8_L1_N14_7= 30'h3ffb99c2,  w8_L1_N14_8= 30'h3ff86738,  w8_L1_N14_9= 30'h3ffb028e,  w8_L1_N14_10= 30'h3ffb36c6,  w8_L1_N14_11= 30'h3ffad595,  w8_L1_N14_12= 30'h3ffc69e8,  w8_L1_N14_13= 30'h3ffb881e,  w8_L1_N14_14= 30'h3ffbf946,  w8_L1_N14_15= 30'h3ffb9cf7,  w8_L1_N14_16= 30'h3ffb0316;
reg [29:0] w8_L1_N15_0= 30'h00026e47,  w8_L1_N15_1= 30'h00013aa2,  w8_L1_N15_2= 30'h000170ae,  w8_L1_N15_3= 30'h3ffbb302,  w8_L1_N15_4= 30'h3ff94b10,  w8_L1_N15_5= 30'h3ffcadad,  w8_L1_N15_6= 30'h3ff84d34,  w8_L1_N15_7= 30'h3ff95f60,  w8_L1_N15_8= 30'h3ffa611a,  w8_L1_N15_9= 30'h3ff8b6f4,  w8_L1_N15_10= 30'h3ffbb92a,  w8_L1_N15_11= 30'h3ff8f062,  w8_L1_N15_12= 30'h3ffc8e73,  w8_L1_N15_13= 30'h3ff9fb8a,  w8_L1_N15_14= 30'h3ffcab21,  w8_L1_N15_15= 30'h3ff9ea89,  w8_L1_N15_16= 30'h3ff93fae;
reg [29:0] w8_L1_N16_0= 30'h00000000,  w8_L1_N16_1= 30'h00000000,  w8_L1_N16_2= 30'h00000000,  w8_L1_N16_3= 30'h00000000,  w8_L1_N16_4= 30'h00000000,  w8_L1_N16_5= 30'h00000000,  w8_L1_N16_6= 30'h00000000,  w8_L1_N16_7= 30'h00000000,  w8_L1_N16_8= 30'h00000000,  w8_L1_N16_9= 30'h00000000,  w8_L1_N16_10= 30'h00000000,  w8_L1_N16_11= 30'h00000000,  w8_L1_N16_12= 30'h00000000,  w8_L1_N16_13= 30'h00000000,  w8_L1_N16_14= 30'h00000000,  w8_L1_N16_15= 30'h00000000,  w8_L1_N16_16= 30'h00000000;
reg [29:0] w8_L1_N17_0= 30'h00000000,  w8_L1_N17_1= 30'h000062be,  w8_L1_N17_2= 30'h00000000,  w8_L1_N17_3= 30'h00000000,  w8_L1_N17_4= 30'h00000000,  w8_L1_N17_5= 30'h00000000,  w8_L1_N17_6= 30'h00000000,  w8_L1_N17_7= 30'h00000000,  w8_L1_N17_8= 30'h00000000,  w8_L1_N17_9= 30'h00000000,  w8_L1_N17_10= 30'h00000000,  w8_L1_N17_11= 30'h00000000,  w8_L1_N17_12= 30'h00000000,  w8_L1_N17_13= 30'h00000000,  w8_L1_N17_14= 30'h00000000,  w8_L1_N17_15= 30'h00000000,  w8_L1_N17_16= 30'h00000000;
reg [29:0] w8_L1_N18_0= 30'h00000000,  w8_L1_N18_1= 30'h00000000,  w8_L1_N18_2= 30'h00000000,  w8_L1_N18_3= 30'h00000000,  w8_L1_N18_4= 30'h00000000,  w8_L1_N18_5= 30'h00000000,  w8_L1_N18_6= 30'h00000000,  w8_L1_N18_7= 30'h00000000,  w8_L1_N18_8= 30'h00000000,  w8_L1_N18_9= 30'h00000000,  w8_L1_N18_10= 30'h00000000,  w8_L1_N18_11= 30'h00000000,  w8_L1_N18_12= 30'h00000000,  w8_L1_N18_13= 30'h00000000,  w8_L1_N18_14= 30'h00000000,  w8_L1_N18_15= 30'h00000000,  w8_L1_N18_16= 30'h00000000;
reg [29:0] w8_L1_N19_0= 30'h3ffb9d86,  w8_L1_N19_1= 30'h3fff7de1,  w8_L1_N19_2= 30'h000039a6,  w8_L1_N19_3= 30'h000c9405,  w8_L1_N19_4= 30'h000f44d9,  w8_L1_N19_5= 30'h000a56de,  w8_L1_N19_6= 30'h0010d3b2,  w8_L1_N19_7= 30'h000f366d,  w8_L1_N19_8= 30'h000f62a3,  w8_L1_N19_9= 30'h001088e8,  w8_L1_N19_10= 30'h000c9131,  w8_L1_N19_11= 30'h001040ec,  w8_L1_N19_12= 30'h000a5c40,  w8_L1_N19_13= 30'h000f62c1,  w8_L1_N19_14= 30'h000a21ab,  w8_L1_N19_15= 30'h000dcbc4,  w8_L1_N19_16= 30'h000f520b;
reg [29:0] w8_L1_N20_0= 30'h00054e31,  w8_L1_N20_1= 30'h0004ec40,  w8_L1_N20_2= 30'h3fff36a0,  w8_L1_N20_3= 30'h3fe661e0,  w8_L1_N20_4= 30'h3fe4455b,  w8_L1_N20_5= 30'h3fe8eb2d,  w8_L1_N20_6= 30'h3fdeb97d,  w8_L1_N20_7= 30'h3fe5f851,  w8_L1_N20_8= 30'h3fe23204,  w8_L1_N20_9= 30'h3fe473d4,  w8_L1_N20_10= 30'h3fe63080,  w8_L1_N20_11= 30'h3fe5ecf9,  w8_L1_N20_12= 30'h3fe8f5d0,  w8_L1_N20_13= 30'h3fe58661,  w8_L1_N20_14= 30'h3fe82e73,  w8_L1_N20_15= 30'h3fe5cfcd,  w8_L1_N20_16= 30'h3fe5a778;
reg [29:0] w8_L1_N21_0= 30'h3ffe15c8,  w8_L1_N21_1= 30'h00012f78,  w8_L1_N21_2= 30'h3fffd708,  w8_L1_N21_3= 30'h0013e97b,  w8_L1_N21_4= 30'h0015df8a,  w8_L1_N21_5= 30'h0010c5de,  w8_L1_N21_6= 30'h00180bff,  w8_L1_N21_7= 30'h0014b20d,  w8_L1_N21_8= 30'h001621a8,  w8_L1_N21_9= 30'h001728e9,  w8_L1_N21_10= 30'h0013ea33,  w8_L1_N21_11= 30'h0016bc80,  w8_L1_N21_12= 30'h0011309d,  w8_L1_N21_13= 30'h00144d9b,  w8_L1_N21_14= 30'h0012441a,  w8_L1_N21_15= 30'h0016189d,  w8_L1_N21_16= 30'h001605fb;
reg [29:0] w8_L1_N22_0= 30'h3ffc172f,  w8_L1_N22_1= 30'h0000492a,  w8_L1_N22_2= 30'h3ffdfe43,  w8_L1_N22_3= 30'h001a2e1e,  w8_L1_N22_4= 30'h001d5458,  w8_L1_N22_5= 30'h001964c0,  w8_L1_N22_6= 30'h0021d54b,  w8_L1_N22_7= 30'h001a89d7,  w8_L1_N22_8= 30'h001e3400,  w8_L1_N22_9= 30'h001d0c22,  w8_L1_N22_10= 30'h001b24a7,  w8_L1_N22_11= 30'h001c1872,  w8_L1_N22_12= 30'h0018a39c,  w8_L1_N22_13= 30'h001aa22d,  w8_L1_N22_14= 30'h0018e870,  w8_L1_N22_15= 30'h001b3fa8,  w8_L1_N22_16= 30'h001d5c7f;
reg [29:0] w8_L1_N23_0= 30'h00000000,  w8_L1_N23_1= 30'h00000000,  w8_L1_N23_2= 30'h00000000,  w8_L1_N23_3= 30'h00000000,  w8_L1_N23_4= 30'h00000000,  w8_L1_N23_5= 30'h00000000,  w8_L1_N23_6= 30'h00000000,  w8_L1_N23_7= 30'h00000000,  w8_L1_N23_8= 30'h00000000,  w8_L1_N23_9= 30'h00000000,  w8_L1_N23_10= 30'h00000000,  w8_L1_N23_11= 30'h00000000,  w8_L1_N23_12= 30'h00000000,  w8_L1_N23_13= 30'h00000000,  w8_L1_N23_14= 30'h00000000,  w8_L1_N23_15= 30'h00000000,  w8_L1_N23_16= 30'h00000000;
reg [29:0] w8_L1_N24_0= 30'h00000000,  w8_L1_N24_1= 30'h00000000,  w8_L1_N24_2= 30'h00000000,  w8_L1_N24_3= 30'h00000000,  w8_L1_N24_4= 30'h00000000,  w8_L1_N24_5= 30'h00000000,  w8_L1_N24_6= 30'h00000000,  w8_L1_N24_7= 30'h00000000,  w8_L1_N24_8= 30'h00000000,  w8_L1_N24_9= 30'h00000000,  w8_L1_N24_10= 30'h00000000,  w8_L1_N24_11= 30'h00000000,  w8_L1_N24_12= 30'h00000000,  w8_L1_N24_13= 30'h00000000,  w8_L1_N24_14= 30'h00000000,  w8_L1_N24_15= 30'h00000000,  w8_L1_N24_16= 30'h00000000;
reg [29:0] w8_L1_N25_0= 30'h3ffa6a5a,  w8_L1_N25_1= 30'h3fff1e83,  w8_L1_N25_2= 30'h3fff6a6a,  w8_L1_N25_3= 30'h00194444,  w8_L1_N25_4= 30'h001af554,  w8_L1_N25_5= 30'h0018c1b5,  w8_L1_N25_6= 30'h00221e3e,  w8_L1_N25_7= 30'h001a71c7,  w8_L1_N25_8= 30'h001e5470,  w8_L1_N25_9= 30'h001b23ce,  w8_L1_N25_10= 30'h0018c951,  w8_L1_N25_11= 30'h001bc32a,  w8_L1_N25_12= 30'h00181f01,  w8_L1_N25_13= 30'h001a6b26,  w8_L1_N25_14= 30'h0018c3eb,  w8_L1_N25_15= 30'h001af74e,  w8_L1_N25_16= 30'h001b175d;
reg [29:0] w8_L1_N26_0= 30'h0002a408,  w8_L1_N26_1= 30'h0003c584,  w8_L1_N26_2= 30'h3fff1dcf,  w8_L1_N26_3= 30'h3ffe41d7,  w8_L1_N26_4= 30'h3ffce3d5,  w8_L1_N26_5= 30'h3ffecb17,  w8_L1_N26_6= 30'h3ffb5eae,  w8_L1_N26_7= 30'h3ffd6af3,  w8_L1_N26_8= 30'h3ffd4157,  w8_L1_N26_9= 30'h3ffd043a,  w8_L1_N26_10= 30'h3ffe412b,  w8_L1_N26_11= 30'h3ffce2de,  w8_L1_N26_12= 30'h3ffee9fe,  w8_L1_N26_13= 30'h3ffd87bf,  w8_L1_N26_14= 30'h3ffec9eb,  w8_L1_N26_15= 30'h3ffd6737,  w8_L1_N26_16= 30'h3ffcf6e6;
reg [29:0] w8_L1_N27_0= 30'h3ff7ce2b,  w8_L1_N27_1= 30'h0005db36,  w8_L1_N27_2= 30'h3ffe7f29,  w8_L1_N27_3= 30'h00174843,  w8_L1_N27_4= 30'h001a4111,  w8_L1_N27_5= 30'h00175251,  w8_L1_N27_6= 30'h001c47e0,  w8_L1_N27_7= 30'h001c482d,  w8_L1_N27_8= 30'h001f09bb,  w8_L1_N27_9= 30'h001a6dfc,  w8_L1_N27_10= 30'h0015e1fa,  w8_L1_N27_11= 30'h001a2a90,  w8_L1_N27_12= 30'h001625aa,  w8_L1_N27_13= 30'h0018e434,  w8_L1_N27_14= 30'h00178949,  w8_L1_N27_15= 30'h001b6111,  w8_L1_N27_16= 30'h001bbcf8;
reg [29:0] w8_L1_N28_0= 30'h0005aaba,  w8_L1_N28_1= 30'h00005945,  w8_L1_N28_2= 30'h0001e0b4,  w8_L1_N28_3= 30'h3ffe5a6b,  w8_L1_N28_4= 30'h3ffcef3f,  w8_L1_N28_5= 30'h3ffeba0a,  w8_L1_N28_6= 30'h3ffbae61,  w8_L1_N28_7= 30'h3ffd4bbb,  w8_L1_N28_8= 30'h3ffd4a03,  w8_L1_N28_9= 30'h3ffcfcd9,  w8_L1_N28_10= 30'h3ffe5899,  w8_L1_N28_11= 30'h3ffcef6a,  w8_L1_N28_12= 30'h3ffee1e2,  w8_L1_N28_13= 30'h3ffd5386,  w8_L1_N28_14= 30'h3ffebb01,  w8_L1_N28_15= 30'h3ffd56aa,  w8_L1_N28_16= 30'h3ffd1667;
reg [29:0] w8_L1_N29_0= 30'h3ffb7c5b,  w8_L1_N29_1= 30'h00011d1c,  w8_L1_N29_2= 30'h3ffddee1,  w8_L1_N29_3= 30'h0014df09,  w8_L1_N29_4= 30'h00167630,  w8_L1_N29_5= 30'h00148c36,  w8_L1_N29_6= 30'h001d6489,  w8_L1_N29_7= 30'h00183b90,  w8_L1_N29_8= 30'h001a81b9,  w8_L1_N29_9= 30'h0018246a,  w8_L1_N29_10= 30'h00151caa,  w8_L1_N29_11= 30'h0019245f,  w8_L1_N29_12= 30'h0013ef45,  w8_L1_N29_13= 30'h0016da45,  w8_L1_N29_14= 30'h00135963,  w8_L1_N29_15= 30'h0017d249,  w8_L1_N29_16= 30'h00199e4f;
reg [29:0] w8_L1_N30_0= 30'h00035e23,  w8_L1_N30_1= 30'h000198e7,  w8_L1_N30_2= 30'h3ffe8b61,  w8_L1_N30_3= 30'h3fe805fd,  w8_L1_N30_4= 30'h3fe627e5,  w8_L1_N30_5= 30'h3feaf748,  w8_L1_N30_6= 30'h3fe11a80,  w8_L1_N30_7= 30'h3fe77f85,  w8_L1_N30_8= 30'h3fe27250,  w8_L1_N30_9= 30'h3fe561b1,  w8_L1_N30_10= 30'h3fe6e038,  w8_L1_N30_11= 30'h3fe4cec7,  w8_L1_N30_12= 30'h3fea22b8,  w8_L1_N30_13= 30'h3fe5e345,  w8_L1_N30_14= 30'h3fea6b6c,  w8_L1_N30_15= 30'h3fe7bbe5,  w8_L1_N30_16= 30'h3fe46870;
reg [29:0] w8_L1_N31_0= 30'h00000000,  w8_L1_N31_1= 30'h00000000,  w8_L1_N31_2= 30'h00000000,  w8_L1_N31_3= 30'h00000000,  w8_L1_N31_4= 30'h00000000,  w8_L1_N31_5= 30'h00000000,  w8_L1_N31_6= 30'h00000000,  w8_L1_N31_7= 30'h00000000,  w8_L1_N31_8= 30'h00000000,  w8_L1_N31_9= 30'h00000000,  w8_L1_N31_10= 30'h00000000,  w8_L1_N31_11= 30'h00000000,  w8_L1_N31_12= 30'h00000000,  w8_L1_N31_13= 30'h00000000,  w8_L1_N31_14= 30'h00000000,  w8_L1_N31_15= 30'h00000000,  w8_L1_N31_16= 30'h00000000;
reg [29:0] w8_L1_N32_0= 30'h3ffb9888,  w8_L1_N32_1= 30'h3ffcae1d,  w8_L1_N32_2= 30'h00026972,  w8_L1_N32_3= 30'h000625c6,  w8_L1_N32_4= 30'h0009967b,  w8_L1_N32_5= 30'h00058a6c,  w8_L1_N32_6= 30'h000b19af,  w8_L1_N32_7= 30'h00082306,  w8_L1_N32_8= 30'h00088efd,  w8_L1_N32_9= 30'h00097fdd,  w8_L1_N32_10= 30'h0006471d,  w8_L1_N32_11= 30'h0009dfd2,  w8_L1_N32_12= 30'h0005417c,  w8_L1_N32_13= 30'h00097e99,  w8_L1_N32_14= 30'h0005abc9,  w8_L1_N32_15= 30'h00089fb3,  w8_L1_N32_16= 30'h000997dd;
reg [29:0] w8_L1_N33_0= 30'h0000f225,  w8_L1_N33_1= 30'h0000c65a,  w8_L1_N33_2= 30'h3ffe3942,  w8_L1_N33_3= 30'h001c9782,  w8_L1_N33_4= 30'h001cbd34,  w8_L1_N33_5= 30'h001a95ba,  w8_L1_N33_6= 30'h00235385,  w8_L1_N33_7= 30'h001c6cc4,  w8_L1_N33_8= 30'h0020ca23,  w8_L1_N33_9= 30'h001e32c7,  w8_L1_N33_10= 30'h001c9b90,  w8_L1_N33_11= 30'h001e5aee,  w8_L1_N33_12= 30'h001a4e70,  w8_L1_N33_13= 30'h001c52a7,  w8_L1_N33_14= 30'h001a8551,  w8_L1_N33_15= 30'h001bd75e,  w8_L1_N33_16= 30'h001cf2c6;
reg [29:0] w8_L1_N34_0= 30'h00000000,  w8_L1_N34_1= 30'h00008d8b,  w8_L1_N34_2= 30'h00000000,  w8_L1_N34_3= 30'h00000000,  w8_L1_N34_4= 30'h00000000,  w8_L1_N34_5= 30'h00000000,  w8_L1_N34_6= 30'h00000000,  w8_L1_N34_7= 30'h00000000,  w8_L1_N34_8= 30'h00000000,  w8_L1_N34_9= 30'h00000000,  w8_L1_N34_10= 30'h00000000,  w8_L1_N34_11= 30'h00000000,  w8_L1_N34_12= 30'h00000000,  w8_L1_N34_13= 30'h00000000,  w8_L1_N34_14= 30'h00000000,  w8_L1_N34_15= 30'h00000000,  w8_L1_N34_16= 30'h00000000;
reg [29:0] w8_L1_N35_0= 30'h0001024d,  w8_L1_N35_1= 30'h3ffd8ece,  w8_L1_N35_2= 30'h00016186,  w8_L1_N35_3= 30'h3ff432eb,  w8_L1_N35_4= 30'h3ff0d4f7,  w8_L1_N35_5= 30'h3ff60b94,  w8_L1_N35_6= 30'h3ff0959a,  w8_L1_N35_7= 30'h3ff1e2aa,  w8_L1_N35_8= 30'h3ff1b058,  w8_L1_N35_9= 30'h3ff06560,  w8_L1_N35_10= 30'h3ff463fb,  w8_L1_N35_11= 30'h3ff1685d,  w8_L1_N35_12= 30'h3ff4d3be,  w8_L1_N35_13= 30'h3ff24c34,  w8_L1_N35_14= 30'h3ff67856,  w8_L1_N35_15= 30'h3ff22d28,  w8_L1_N35_16= 30'h3ff02e5d;
reg [29:0] w8_L1_N36_0= 30'h3ffdc9f4,  w8_L1_N36_1= 30'h3ffe76fb,  w8_L1_N36_2= 30'h00035cc4,  w8_L1_N36_3= 30'h3ff764c5,  w8_L1_N36_4= 30'h3ff3c03d,  w8_L1_N36_5= 30'h3ff8fa4d,  w8_L1_N36_6= 30'h3ff437f8,  w8_L1_N36_7= 30'h3ff4b9fe,  w8_L1_N36_8= 30'h3ff56923,  w8_L1_N36_9= 30'h3ff3a93d,  w8_L1_N36_10= 30'h3ff78c5d,  w8_L1_N36_11= 30'h3ff3b508,  w8_L1_N36_12= 30'h3ff81b8c,  w8_L1_N36_13= 30'h3ff5dc58,  w8_L1_N36_14= 30'h3ff8cda7,  w8_L1_N36_15= 30'h3ff4b814,  w8_L1_N36_16= 30'h3ff3fd6e;
reg [29:0] w8_L1_N37_0= 30'h00000000,  w8_L1_N37_1= 30'h00012e7f,  w8_L1_N37_2= 30'h00000000,  w8_L1_N37_3= 30'h00000000,  w8_L1_N37_4= 30'h00000000,  w8_L1_N37_5= 30'h00000000,  w8_L1_N37_6= 30'h00000000,  w8_L1_N37_7= 30'h00000000,  w8_L1_N37_8= 30'h00000000,  w8_L1_N37_9= 30'h00000000,  w8_L1_N37_10= 30'h00000000,  w8_L1_N37_11= 30'h00000000,  w8_L1_N37_12= 30'h00000000,  w8_L1_N37_13= 30'h00000000,  w8_L1_N37_14= 30'h00000000,  w8_L1_N37_15= 30'h00000000,  w8_L1_N37_16= 30'h00000000;
reg [29:0] w8_L1_N38_0= 30'h00000000,  w8_L1_N38_1= 30'h00000000,  w8_L1_N38_2= 30'h00000000,  w8_L1_N38_3= 30'h00000000,  w8_L1_N38_4= 30'h00000000,  w8_L1_N38_5= 30'h00000000,  w8_L1_N38_6= 30'h00000000,  w8_L1_N38_7= 30'h00000000,  w8_L1_N38_8= 30'h00000000,  w8_L1_N38_9= 30'h00000000,  w8_L1_N38_10= 30'h00000000,  w8_L1_N38_11= 30'h00000000,  w8_L1_N38_12= 30'h00000000,  w8_L1_N38_13= 30'h00000000,  w8_L1_N38_14= 30'h00000000,  w8_L1_N38_15= 30'h00000000,  w8_L1_N38_16= 30'h00000000;
reg [29:0] w8_L1_N39_0= 30'h0000f098,  w8_L1_N39_1= 30'h00025984,  w8_L1_N39_2= 30'h0003ac9e,  w8_L1_N39_3= 30'h3ff6092f,  w8_L1_N39_4= 30'h3ff2afe6,  w8_L1_N39_5= 30'h3ff78f8c,  w8_L1_N39_6= 30'h3ff23f20,  w8_L1_N39_7= 30'h3ff340c3,  w8_L1_N39_8= 30'h3ff395c9,  w8_L1_N39_9= 30'h3ff2a1ba,  w8_L1_N39_10= 30'h3ff5e2f5,  w8_L1_N39_11= 30'h3ff323e0,  w8_L1_N39_12= 30'h3ff67c98,  w8_L1_N39_13= 30'h3ff3671f,  w8_L1_N39_14= 30'h3ff7c905,  w8_L1_N39_15= 30'h3ff3ea65,  w8_L1_N39_16= 30'h3ff1dc12;
reg [29:0] w8_L1_N40_0= 30'h3ff82ec1,  w8_L1_N40_1= 30'h000165a1,  w8_L1_N40_2= 30'h0000980e,  w8_L1_N40_3= 30'h00150877,  w8_L1_N40_4= 30'h0016f3e8,  w8_L1_N40_5= 30'h00135bc2,  w8_L1_N40_6= 30'h001e2d5f,  w8_L1_N40_7= 30'h00188886,  w8_L1_N40_8= 30'h0019bd6e,  w8_L1_N40_9= 30'h00183da8,  w8_L1_N40_10= 30'h00131303,  w8_L1_N40_11= 30'h00181f78,  w8_L1_N40_12= 30'h0011b0a6,  w8_L1_N40_13= 30'h0016b6be,  w8_L1_N40_14= 30'h00144cbf,  w8_L1_N40_15= 30'h0017eebc,  w8_L1_N40_16= 30'h0018f24b;
reg [29:0] w8_L1_N41_0= 30'h3ffae15b,  w8_L1_N41_1= 30'h000029c5,  w8_L1_N41_2= 30'h0002de1c,  w8_L1_N41_3= 30'h00076347,  w8_L1_N41_4= 30'h000b5696,  w8_L1_N41_5= 30'h0006e7bb,  w8_L1_N41_6= 30'h000cbfdc,  w8_L1_N41_7= 30'h000aeb23,  w8_L1_N41_8= 30'h000a42b7,  w8_L1_N41_9= 30'h000b3cf1,  w8_L1_N41_10= 30'h0007b2a3,  w8_L1_N41_11= 30'h000a8a42,  w8_L1_N41_12= 30'h0007294e,  w8_L1_N41_13= 30'h000b0b6c,  w8_L1_N41_14= 30'h00066d09,  w8_L1_N41_15= 30'h000a5035,  w8_L1_N41_16= 30'h000a966a;
reg [29:0] w8_L1_N42_0= 30'h00010cb4,  w8_L1_N42_1= 30'h00000688,  w8_L1_N42_2= 30'h0003e414,  w8_L1_N42_3= 30'h3ff875aa,  w8_L1_N42_4= 30'h3ff52807,  w8_L1_N42_5= 30'h3ffa20fa,  w8_L1_N42_6= 30'h3ff6234a,  w8_L1_N42_7= 30'h3ff5dc2d,  w8_L1_N42_8= 30'h3ff6cbdc,  w8_L1_N42_9= 30'h3ff5b105,  w8_L1_N42_10= 30'h3ff895f1,  w8_L1_N42_11= 30'h3ff5bde7,  w8_L1_N42_12= 30'h3ff93a0b,  w8_L1_N42_13= 30'h3ff6c0e6,  w8_L1_N42_14= 30'h3ffa26f4,  w8_L1_N42_15= 30'h3ff60830,  w8_L1_N42_16= 30'h3ff4ea5d;
reg [29:0] w8_L1_N43_0= 30'h000063f7,  w8_L1_N43_1= 30'h000142a6,  w8_L1_N43_2= 30'h3ffffd52,  w8_L1_N43_3= 30'h000ac6d8,  w8_L1_N43_4= 30'h000d0c70,  w8_L1_N43_5= 30'h0008e566,  w8_L1_N43_6= 30'h000dec70,  w8_L1_N43_7= 30'h000cb927,  w8_L1_N43_8= 30'h000d1e63,  w8_L1_N43_9= 30'h000ea4f6,  w8_L1_N43_10= 30'h000a8fd4,  w8_L1_N43_11= 30'h000cde46,  w8_L1_N43_12= 30'h0009c845,  w8_L1_N43_13= 30'h000c8fdf,  w8_L1_N43_14= 30'h0009327f,  w8_L1_N43_15= 30'h000da66e,  w8_L1_N43_16= 30'h000d5bd3;
reg [29:0] w8_L1_N44_0= 30'h3fffc40c,  w8_L1_N44_1= 30'h3fffae78,  w8_L1_N44_2= 30'h0002a6dc,  w8_L1_N44_3= 30'h3ff9221f,  w8_L1_N44_4= 30'h3ff6833f,  w8_L1_N44_5= 30'h3ffa95b2,  w8_L1_N44_6= 30'h3ff7660a,  w8_L1_N44_7= 30'h3ff7d8c7,  w8_L1_N44_8= 30'h3ff7976a,  w8_L1_N44_9= 30'h3ff69fad,  w8_L1_N44_10= 30'h3ff90129,  w8_L1_N44_11= 30'h3ff6e135,  w8_L1_N44_12= 30'h3ff9bc4c,  w8_L1_N44_13= 30'h3ff76e52,  w8_L1_N44_14= 30'h3ffa8dac,  w8_L1_N44_15= 30'h3ff6ece6,  w8_L1_N44_16= 30'h3ff641d4;
reg [29:0] w8_L1_N45_0= 30'h00025b35,  w8_L1_N45_1= 30'h00054988,  w8_L1_N45_2= 30'h3fffe9f9,  w8_L1_N45_3= 30'h3fe5c93d,  w8_L1_N45_4= 30'h3fe50f03,  w8_L1_N45_5= 30'h3fe84bd9,  w8_L1_N45_6= 30'h3fdf31ad,  w8_L1_N45_7= 30'h3fe4503e,  w8_L1_N45_8= 30'h3fe214c7,  w8_L1_N45_9= 30'h3fe3b996,  w8_L1_N45_10= 30'h3fe5d968,  w8_L1_N45_11= 30'h3fe5d8a4,  w8_L1_N45_12= 30'h3fe7e3db,  w8_L1_N45_13= 30'h3fe48c37,  w8_L1_N45_14= 30'h3fe6a78c,  w8_L1_N45_15= 30'h3fe4f830,  w8_L1_N45_16= 30'h3fe402fa;
reg [29:0] w8_L1_N46_0= 30'h3ffff4fb,  w8_L1_N46_1= 30'h3ffeb70e,  w8_L1_N46_2= 30'h0000c4b0,  w8_L1_N46_3= 30'h0010b382,  w8_L1_N46_4= 30'h0013d072,  w8_L1_N46_5= 30'h000d6409,  w8_L1_N46_6= 30'h001534a5,  w8_L1_N46_7= 30'h00114265,  w8_L1_N46_8= 30'h0012e858,  w8_L1_N46_9= 30'h0013754a,  w8_L1_N46_10= 30'h0010ca5e,  w8_L1_N46_11= 30'h001417dc,  w8_L1_N46_12= 30'h000ef320,  w8_L1_N46_13= 30'h0012c421,  w8_L1_N46_14= 30'h000d75b9,  w8_L1_N46_15= 30'h0012422f,  w8_L1_N46_16= 30'h0012a245;
reg [29:0] w8_L1_N47_0= 30'h3ffa98c7,  w8_L1_N47_1= 30'h00019dc1,  w8_L1_N47_2= 30'h3ffe8b4b,  w8_L1_N47_3= 30'h00125559,  w8_L1_N47_4= 30'h001553e3,  w8_L1_N47_5= 30'h0010b7fb,  w8_L1_N47_6= 30'h001833b6,  w8_L1_N47_7= 30'h0014402d,  w8_L1_N47_8= 30'h0015f934,  w8_L1_N47_9= 30'h0014a1cb,  w8_L1_N47_10= 30'h0011fe00,  w8_L1_N47_11= 30'h0015707f,  w8_L1_N47_12= 30'h0010eaf6,  w8_L1_N47_13= 30'h00159a21,  w8_L1_N47_14= 30'h00105504,  w8_L1_N47_15= 30'h0013c995,  w8_L1_N47_16= 30'h00161b18;
reg [29:0] w8_L1_N48_0= 30'h00038fbc,  w8_L1_N48_1= 30'h000282a2,  w8_L1_N48_2= 30'h3fff7d76,  w8_L1_N48_3= 30'h3ffdef72,  w8_L1_N48_4= 30'h3ffc4c38,  w8_L1_N48_5= 30'h3ffe57ca,  w8_L1_N48_6= 30'h3ffa667a,  w8_L1_N48_7= 30'h3ffcd100,  w8_L1_N48_8= 30'h3ffc7f05,  w8_L1_N48_9= 30'h3ffc6031,  w8_L1_N48_10= 30'h3ffdf465,  w8_L1_N48_11= 30'h3ffc4bc2,  w8_L1_N48_12= 30'h3ffe9aa7,  w8_L1_N48_13= 30'h3ffcabe3,  w8_L1_N48_14= 30'h3ffe5b2d,  w8_L1_N48_15= 30'h3ffca85f,  w8_L1_N48_16= 30'h3ffc6a34;
reg [29:0] w8_L1_N49_0= 30'h00000000,  w8_L1_N49_1= 30'h000108f0,  w8_L1_N49_2= 30'h00000000,  w8_L1_N49_3= 30'h00000000,  w8_L1_N49_4= 30'h00000000,  w8_L1_N49_5= 30'h00000000,  w8_L1_N49_6= 30'h00000000,  w8_L1_N49_7= 30'h00000000,  w8_L1_N49_8= 30'h00000000,  w8_L1_N49_9= 30'h00000000,  w8_L1_N49_10= 30'h00000000,  w8_L1_N49_11= 30'h00000000,  w8_L1_N49_12= 30'h00000000,  w8_L1_N49_13= 30'h00000000,  w8_L1_N49_14= 30'h00000000,  w8_L1_N49_15= 30'h00000000,  w8_L1_N49_16= 30'h00000000;
reg [29:0] w8_L1_N50_0= 30'h000529ff,  w8_L1_N50_1= 30'h0002b4e4,  w8_L1_N50_2= 30'h3ffdecc8,  w8_L1_N50_3= 30'h00199447,  w8_L1_N50_4= 30'h001bbc57,  w8_L1_N50_5= 30'h0017da81,  w8_L1_N50_6= 30'h002190a8,  w8_L1_N50_7= 30'h001af325,  w8_L1_N50_8= 30'h001eba02,  w8_L1_N50_9= 30'h001c90e1,  w8_L1_N50_10= 30'h00199c58,  w8_L1_N50_11= 30'h001c1dad,  w8_L1_N50_12= 30'h00181b9d,  w8_L1_N50_13= 30'h001a4f76,  w8_L1_N50_14= 30'h001808d1,  w8_L1_N50_15= 30'h001afe07,  w8_L1_N50_16= 30'h001cb62a;
reg [29:0] w8_L1_N51_0= 30'h00000000,  w8_L1_N51_1= 30'h00000000,  w8_L1_N51_2= 30'h00000000,  w8_L1_N51_3= 30'h00000000,  w8_L1_N51_4= 30'h00000000,  w8_L1_N51_5= 30'h00000000,  w8_L1_N51_6= 30'h00000000,  w8_L1_N51_7= 30'h00000000,  w8_L1_N51_8= 30'h00000000,  w8_L1_N51_9= 30'h00000000,  w8_L1_N51_10= 30'h00000000,  w8_L1_N51_11= 30'h00000000,  w8_L1_N51_12= 30'h00000000,  w8_L1_N51_13= 30'h00000000,  w8_L1_N51_14= 30'h00000000,  w8_L1_N51_15= 30'h00000000,  w8_L1_N51_16= 30'h00000000;
reg [29:0] w8_L1_N52_0= 30'h00044c32,  w8_L1_N52_1= 30'h000310d2,  w8_L1_N52_2= 30'h3ffe3520,  w8_L1_N52_3= 30'h3fe61d3e,  w8_L1_N52_4= 30'h3fe43572,  w8_L1_N52_5= 30'h3fe61254,  w8_L1_N52_6= 30'h3fdc59bc,  w8_L1_N52_7= 30'h3fe38667,  w8_L1_N52_8= 30'h3fe12d49,  w8_L1_N52_9= 30'h3fe494d0,  w8_L1_N52_10= 30'h3fe64330,  w8_L1_N52_11= 30'h3fe483b7,  w8_L1_N52_12= 30'h3fe72069,  w8_L1_N52_13= 30'h3fe66ef8,  w8_L1_N52_14= 30'h3fe627bb,  w8_L1_N52_15= 30'h3fe39be4,  w8_L1_N52_16= 30'h3fe28787;
reg [29:0] w8_L1_N53_0= 30'h0007f09f,  w8_L1_N53_1= 30'h00057e85,  w8_L1_N53_2= 30'h3ffec6bd,  w8_L1_N53_3= 30'h000cde0e,  w8_L1_N53_4= 30'h000e6412,  w8_L1_N53_5= 30'h000b00c8,  w8_L1_N53_6= 30'h0011b679,  w8_L1_N53_7= 30'h000d50cc,  w8_L1_N53_8= 30'h0010764f,  w8_L1_N53_9= 30'h000ee8ae,  w8_L1_N53_10= 30'h000cde9c,  w8_L1_N53_11= 30'h000e6427,  w8_L1_N53_12= 30'h000b84ab,  w8_L1_N53_13= 30'h000cf97d,  w8_L1_N53_14= 30'h000b00c8,  w8_L1_N53_15= 30'h000d50ce,  w8_L1_N53_16= 30'h000ee8b1;
reg [29:0] w8_L1_N54_0= 30'h0003fb13,  w8_L1_N54_1= 30'h0000dbf0,  w8_L1_N54_2= 30'h0002ec03,  w8_L1_N54_3= 30'h3ffa2fd7,  w8_L1_N54_4= 30'h3ff6af89,  w8_L1_N54_5= 30'h3ffb1d6d,  w8_L1_N54_6= 30'h3ff6a0ec,  w8_L1_N54_7= 30'h3ff7c58e,  w8_L1_N54_8= 30'h3ff86b0c,  w8_L1_N54_9= 30'h3ff6b14d,  w8_L1_N54_10= 30'h3ffa1994,  w8_L1_N54_11= 30'h3ff6aa8b,  w8_L1_N54_12= 30'h3ffac390,  w8_L1_N54_13= 30'h3ff7ec4c,  w8_L1_N54_14= 30'h3ffb3b28,  w8_L1_N54_15= 30'h3ff7bdc7,  w8_L1_N54_16= 30'h3ff68b63;
reg [29:0] w8_L1_N55_0= 30'h3ffcc92d,  w8_L1_N55_1= 30'h3ffe64c2,  w8_L1_N55_2= 30'h0001ceaa,  w8_L1_N55_3= 30'h0004b521,  w8_L1_N55_4= 30'h000767b0,  w8_L1_N55_5= 30'h0003dc36,  w8_L1_N55_6= 30'h0007e03e,  w8_L1_N55_7= 30'h0006c2ae,  w8_L1_N55_8= 30'h0006c709,  w8_L1_N55_9= 30'h000771d8,  w8_L1_N55_10= 30'h00049323,  w8_L1_N55_11= 30'h0006e5d0,  w8_L1_N55_12= 30'h00040ec9,  w8_L1_N55_13= 30'h0006fed4,  w8_L1_N55_14= 30'h0003ebd2,  w8_L1_N55_15= 30'h00068268,  w8_L1_N55_16= 30'h00078e04;
reg [29:0] w8_L1_N56_0= 30'h00057a5b,  w8_L1_N56_1= 30'h000141b4,  w8_L1_N56_2= 30'h3ffe8f3a,  w8_L1_N56_3= 30'h001b6658,  w8_L1_N56_4= 30'h001d6850,  w8_L1_N56_5= 30'h0019b379,  w8_L1_N56_6= 30'h0023396f,  w8_L1_N56_7= 30'h001bfc9a,  w8_L1_N56_8= 30'h0020723b,  w8_L1_N56_9= 30'h001dac4d,  w8_L1_N56_10= 30'h001b11c6,  w8_L1_N56_11= 30'h001d7803,  w8_L1_N56_12= 30'h001a129d,  w8_L1_N56_13= 30'h001ba466,  w8_L1_N56_14= 30'h001a025b,  w8_L1_N56_15= 30'h001c7a6e,  w8_L1_N56_16= 30'h001db0c2;
reg [29:0] w8_L1_N57_0= 30'h00000000,  w8_L1_N57_1= 30'h3fffd209,  w8_L1_N57_2= 30'h3fffe9e4,  w8_L1_N57_3= 30'h00000000,  w8_L1_N57_4= 30'h00000000,  w8_L1_N57_5= 30'h00000000,  w8_L1_N57_6= 30'h00000000,  w8_L1_N57_7= 30'h00000000,  w8_L1_N57_8= 30'h00000000,  w8_L1_N57_9= 30'h00000000,  w8_L1_N57_10= 30'h00000000,  w8_L1_N57_11= 30'h00000000,  w8_L1_N57_12= 30'h00000000,  w8_L1_N57_13= 30'h00000000,  w8_L1_N57_14= 30'h00000000,  w8_L1_N57_15= 30'h00000000,  w8_L1_N57_16= 30'h00000000;
reg [29:0] w8_L1_N58_0= 30'h3ff60653,  w8_L1_N58_1= 30'h0001b47a,  w8_L1_N58_2= 30'h00015e1e,  w8_L1_N58_3= 30'h00146f1f,  w8_L1_N58_4= 30'h0018b120,  w8_L1_N58_5= 30'h0014b7a1,  w8_L1_N58_6= 30'h001ea739,  w8_L1_N58_7= 30'h00171280,  w8_L1_N58_8= 30'h001a96ca,  w8_L1_N58_9= 30'h00181bf2,  w8_L1_N58_10= 30'h0014810d,  w8_L1_N58_11= 30'h0018e208,  w8_L1_N58_12= 30'h00136830,  w8_L1_N58_13= 30'h00159681,  w8_L1_N58_14= 30'h001367f5,  w8_L1_N58_15= 30'h00193014,  w8_L1_N58_16= 30'h0017eb2d;
reg [29:0] w8_L1_N59_0= 30'h3ff6b951,  w8_L1_N59_1= 30'h0006af6d,  w8_L1_N59_2= 30'h3ffeab61,  w8_L1_N59_3= 30'h00173aed,  w8_L1_N59_4= 30'h001cf0c5,  w8_L1_N59_5= 30'h001896b3,  w8_L1_N59_6= 30'h001e9751,  w8_L1_N59_7= 30'h001ef90a,  w8_L1_N59_8= 30'h00208398,  w8_L1_N59_9= 30'h001b3e06,  w8_L1_N59_10= 30'h0018c357,  w8_L1_N59_11= 30'h001b9509,  w8_L1_N59_12= 30'h0018098a,  w8_L1_N59_13= 30'h001b774d,  w8_L1_N59_14= 30'h0019d216,  w8_L1_N59_15= 30'h001e9fe6,  w8_L1_N59_16= 30'h001bf922;
reg [29:0] w8_L1_N60_0= 30'h0000576b,  w8_L1_N60_1= 30'h3ffd90e1,  w8_L1_N60_2= 30'h00002e17,  w8_L1_N60_3= 30'h000f73e6,  w8_L1_N60_4= 30'h001196c2,  w8_L1_N60_5= 30'h000da092,  w8_L1_N60_6= 30'h0015178e,  w8_L1_N60_7= 30'h00113da3,  w8_L1_N60_8= 30'h00138b2c,  w8_L1_N60_9= 30'h0012c4b2,  w8_L1_N60_10= 30'h0010b8d0,  w8_L1_N60_11= 30'h0012115b,  w8_L1_N60_12= 30'h000ea6ec,  w8_L1_N60_13= 30'h0011d5f8,  w8_L1_N60_14= 30'h000d9e5b,  w8_L1_N60_15= 30'h00116fac,  w8_L1_N60_16= 30'h00135c49;

reg [29:0] w8_L2_N1_0= 30'h00000000,  w8_L2_N1_1= 30'h00000000,  w8_L2_N1_2= 30'h00008f4e,  w8_L2_N1_3= 30'h3fff154c,  w8_L2_N1_4= 30'h00000000,  w8_L2_N1_5= 30'h00000000,  w8_L2_N1_6= 30'h00000000,  w8_L2_N1_7= 30'h00007d24,  w8_L2_N1_8= 30'h00008aa1,  w8_L2_N1_9= 30'h3fff5308,  w8_L2_N1_10= 30'h3ffef9bf,  w8_L2_N1_11= 30'h00000000,  w8_L2_N1_12= 30'h0000584c,  w8_L2_N1_13= 30'h00000000,  w8_L2_N1_14= 30'h000006b1,  w8_L2_N1_15= 30'h00000000,  w8_L2_N1_16= 30'h3fffad78,  w8_L2_N1_17= 30'h00000000,  w8_L2_N1_18= 30'h0000f0fb,  w8_L2_N1_19= 30'h00002716,  w8_L2_N1_20= 30'h3fff5162,  w8_L2_N1_21= 30'h000051b8,  w8_L2_N1_22= 30'h00000000,  w8_L2_N1_23= 30'h00000000,  w8_L2_N1_24= 30'h00000000,  w8_L2_N1_25= 30'h3fff0672,  w8_L2_N1_26= 30'h3ffe6b1e,  w8_L2_N1_27= 30'h3fffcfec,  w8_L2_N1_28= 30'h3ffed6c6,  w8_L2_N1_29= 30'h3fff1eae;
reg [29:0] w8_L2_N1_30= 30'h00000000,  w8_L2_N1_31= 30'h3fffe855,  w8_L2_N1_32= 30'h3fffff83,  w8_L2_N1_33= 30'h3fff2d34,  w8_L2_N1_34= 30'h3fffbab4,  w8_L2_N1_35= 30'h3ffff442,  w8_L2_N1_36= 30'h3fffdfdb,  w8_L2_N1_37= 30'h00000000,  w8_L2_N1_38= 30'h3fffa6ab,  w8_L2_N1_39= 30'h00007bcd,  w8_L2_N1_40= 30'h3fff23f0,  w8_L2_N1_41= 30'h3ffe78b4,  w8_L2_N1_42= 30'h00016467,  w8_L2_N1_43= 30'h3ffe7088,  w8_L2_N1_44= 30'h00004564,  w8_L2_N1_45= 30'h00006814,  w8_L2_N1_46= 30'h3fffbb77,  w8_L2_N1_47= 30'h3ffea428,  w8_L2_N1_48= 30'h00000001,  w8_L2_N1_49= 30'h3fff9593,  w8_L2_N1_50= 30'h00000000,  w8_L2_N1_51= 30'h00000000,  w8_L2_N1_52= 30'h00000000,  w8_L2_N1_53= 30'h3ffef437,  w8_L2_N1_54= 30'h0001741d,  w8_L2_N1_55= 30'h3fffe405,  w8_L2_N1_56= 30'h3fffca92,  w8_L2_N1_57= 30'h3fff460f,  w8_L2_N1_58= 30'h0000f89e,  w8_L2_N1_59= 30'h00004f64;
reg [29:0] w8_L2_N2_0= 30'h00000000,  w8_L2_N2_1= 30'h00000000,  w8_L2_N2_2= 30'h00000000,  w8_L2_N2_3= 30'h00000000,  w8_L2_N2_4= 30'h00000000,  w8_L2_N2_5= 30'h00000000,  w8_L2_N2_6= 30'h00000000,  w8_L2_N2_7= 30'h00000000,  w8_L2_N2_8= 30'h00000000,  w8_L2_N2_9= 30'h00000000,  w8_L2_N2_10= 30'h00000000,  w8_L2_N2_11= 30'h00000000,  w8_L2_N2_12= 30'h00000000,  w8_L2_N2_13= 30'h00000000,  w8_L2_N2_14= 30'h00000000,  w8_L2_N2_15= 30'h00000000,  w8_L2_N2_16= 30'h00000000,  w8_L2_N2_17= 30'h00000000,  w8_L2_N2_18= 30'h00000000,  w8_L2_N2_19= 30'h00000000,  w8_L2_N2_20= 30'h00000000,  w8_L2_N2_21= 30'h00000000,  w8_L2_N2_22= 30'h00000000,  w8_L2_N2_23= 30'h00000000,  w8_L2_N2_24= 30'h00000000,  w8_L2_N2_25= 30'h00000000,  w8_L2_N2_26= 30'h00000000,  w8_L2_N2_27= 30'h00000000,  w8_L2_N2_28= 30'h00000000,  w8_L2_N2_29= 30'h00000000;
reg [29:0] w8_L2_N2_30= 30'h00000000,  w8_L2_N2_31= 30'h00000000,  w8_L2_N2_32= 30'h00000000,  w8_L2_N2_33= 30'h00000000,  w8_L2_N2_34= 30'h00000000,  w8_L2_N2_35= 30'h00000000,  w8_L2_N2_36= 30'h00000000,  w8_L2_N2_37= 30'h00000000,  w8_L2_N2_38= 30'h00000000,  w8_L2_N2_39= 30'h00000000,  w8_L2_N2_40= 30'h00000000,  w8_L2_N2_41= 30'h00000000,  w8_L2_N2_42= 30'h00000000,  w8_L2_N2_43= 30'h00000000,  w8_L2_N2_44= 30'h00000000,  w8_L2_N2_45= 30'h00000000,  w8_L2_N2_46= 30'h00000000,  w8_L2_N2_47= 30'h00000000,  w8_L2_N2_48= 30'h00000000,  w8_L2_N2_49= 30'h00000000,  w8_L2_N2_50= 30'h00000000,  w8_L2_N2_51= 30'h00000000,  w8_L2_N2_52= 30'h00000000,  w8_L2_N2_53= 30'h00000000,  w8_L2_N2_54= 30'h00000000,  w8_L2_N2_55= 30'h00000000,  w8_L2_N2_56= 30'h00000000,  w8_L2_N2_57= 30'h00000000,  w8_L2_N2_58= 30'h00000000,  w8_L2_N2_59= 30'h00000000;
reg [29:0] w8_L2_N3_0= 30'h00000000,  w8_L2_N3_1= 30'h00000000,  w8_L2_N3_2= 30'h00028649,  w8_L2_N3_3= 30'h0002e313,  w8_L2_N3_4= 30'h00000000,  w8_L2_N3_5= 30'h00000000,  w8_L2_N3_6= 30'h00000000,  w8_L2_N3_7= 30'h3fff6eae,  w8_L2_N3_8= 30'h000126d9,  w8_L2_N3_9= 30'h3fffdd4d,  w8_L2_N3_10= 30'h3ffe318a,  w8_L2_N3_11= 30'h00000000,  w8_L2_N3_12= 30'h0002e5f8,  w8_L2_N3_13= 30'h00011a92,  w8_L2_N3_14= 30'h0001b3a3,  w8_L2_N3_15= 30'h00000000,  w8_L2_N3_16= 30'h000087e8,  w8_L2_N3_17= 30'h00000000,  w8_L2_N3_18= 30'h3ffe5e6f,  w8_L2_N3_19= 30'h000329ea,  w8_L2_N3_20= 30'h3ffe1da8,  w8_L2_N3_21= 30'h3ffb0a1f,  w8_L2_N3_22= 30'h00000000,  w8_L2_N3_23= 30'h00000000,  w8_L2_N3_24= 30'h3ffbb571,  w8_L2_N3_25= 30'h00012bbf,  w8_L2_N3_26= 30'h3ffb9cd9,  w8_L2_N3_27= 30'h3ffffbac,  w8_L2_N3_28= 30'h3ffe60b3,  w8_L2_N3_29= 30'h0000f669;
reg [29:0] w8_L2_N3_30= 30'h00000000,  w8_L2_N3_31= 30'h0002a3af,  w8_L2_N3_32= 30'h3ff8e58d,  w8_L2_N3_33= 30'h3ffff2ef,  w8_L2_N3_34= 30'h000388d8,  w8_L2_N3_35= 30'h0003a234,  w8_L2_N3_36= 30'h000009e4,  w8_L2_N3_37= 30'h00000000,  w8_L2_N3_38= 30'h0000e2ee,  w8_L2_N3_39= 30'h3ffa585d,  w8_L2_N3_40= 30'h0001e491,  w8_L2_N3_41= 30'h00036da2,  w8_L2_N3_42= 30'h3ffdd68f,  w8_L2_N3_43= 30'h00040315,  w8_L2_N3_44= 30'h00033b69,  w8_L2_N3_45= 30'h3fff77a4,  w8_L2_N3_46= 30'h3fff1834,  w8_L2_N3_47= 30'h00021483,  w8_L2_N3_48= 30'h3fffffe3,  w8_L2_N3_49= 30'h3ffd8876,  w8_L2_N3_50= 30'h00000000,  w8_L2_N3_51= 30'h00028f3d,  w8_L2_N3_52= 30'h3ffc0745,  w8_L2_N3_53= 30'h3fff6f00,  w8_L2_N3_54= 30'h0001b888,  w8_L2_N3_55= 30'h3ff867a9,  w8_L2_N3_56= 30'h00002eb6,  w8_L2_N3_57= 30'h3ffa823b,  w8_L2_N3_58= 30'h3ffadbcb,  w8_L2_N3_59= 30'h3fff5d5d;
reg [29:0] w8_L2_N4_0= 30'h00000000,  w8_L2_N4_1= 30'h00000000,  w8_L2_N4_2= 30'h3fff5463,  w8_L2_N4_3= 30'h3fff2896,  w8_L2_N4_4= 30'h00000000,  w8_L2_N4_5= 30'h00000000,  w8_L2_N4_6= 30'h00000000,  w8_L2_N4_7= 30'h0001f542,  w8_L2_N4_8= 30'h0002179f,  w8_L2_N4_9= 30'h000023b7,  w8_L2_N4_10= 30'h00024022,  w8_L2_N4_11= 30'h00000000,  w8_L2_N4_12= 30'h3fff414e,  w8_L2_N4_13= 30'h000261d9,  w8_L2_N4_14= 30'h3fff9ed8,  w8_L2_N4_15= 30'h00000000,  w8_L2_N4_16= 30'h00000000,  w8_L2_N4_17= 30'h00000000,  w8_L2_N4_18= 30'h00002ac2,  w8_L2_N4_19= 30'h00017337,  w8_L2_N4_20= 30'h000095c8,  w8_L2_N4_21= 30'h0001cef7,  w8_L2_N4_22= 30'h00000000,  w8_L2_N4_23= 30'h00000000,  w8_L2_N4_24= 30'h000053c9,  w8_L2_N4_25= 30'h0000d1ce,  w8_L2_N4_26= 30'h0002edb7,  w8_L2_N4_27= 30'h3fff3dd4,  w8_L2_N4_28= 30'h00022c4f,  w8_L2_N4_29= 30'h00011d46;
reg [29:0] w8_L2_N4_30= 30'h00000000,  w8_L2_N4_31= 30'h3fff4f3c,  w8_L2_N4_32= 30'h000123ce,  w8_L2_N4_33= 30'h00000000,  w8_L2_N4_34= 30'h3fff7343,  w8_L2_N4_35= 30'h3fff7b8c,  w8_L2_N4_36= 30'h00000000,  w8_L2_N4_37= 30'h00000000,  w8_L2_N4_38= 30'h3fff4da9,  w8_L2_N4_39= 30'h00002275,  w8_L2_N4_40= 30'h3fff8cf0,  w8_L2_N4_41= 30'h3fff32cc,  w8_L2_N4_42= 30'h00005bc8,  w8_L2_N4_43= 30'h3fff633a,  w8_L2_N4_44= 30'h0001bddb,  w8_L2_N4_45= 30'h3fff7ae8,  w8_L2_N4_46= 30'h0001d556,  w8_L2_N4_47= 30'h00005453,  w8_L2_N4_48= 30'h00000000,  w8_L2_N4_49= 30'h00014c07,  w8_L2_N4_50= 30'h00000000,  w8_L2_N4_51= 30'h0001b0cf,  w8_L2_N4_52= 30'h00018418,  w8_L2_N4_53= 30'h3fff3d6d,  w8_L2_N4_54= 30'h3fff77f4,  w8_L2_N4_55= 30'h000081fa,  w8_L2_N4_56= 30'h00000000,  w8_L2_N4_57= 30'h3ffff3d8,  w8_L2_N4_58= 30'h000315c4,  w8_L2_N4_59= 30'h3fff71ae;
reg [29:0] w8_L2_N5_0= 30'h00000000,  w8_L2_N5_1= 30'h00000000,  w8_L2_N5_2= 30'h3fffcf9e,  w8_L2_N5_3= 30'h3ffd2b97,  w8_L2_N5_4= 30'h00000000,  w8_L2_N5_5= 30'h00000000,  w8_L2_N5_6= 30'h00000000,  w8_L2_N5_7= 30'h00079785,  w8_L2_N5_8= 30'h3ff0764b,  w8_L2_N5_9= 30'h00005e16,  w8_L2_N5_10= 30'h00075ca1,  w8_L2_N5_11= 30'h00000000,  w8_L2_N5_12= 30'h00006ce7,  w8_L2_N5_13= 30'h3ffc9f1a,  w8_L2_N5_14= 30'h3ffe00aa,  w8_L2_N5_15= 30'h00000000,  w8_L2_N5_16= 30'h00000000,  w8_L2_N5_17= 30'h00000000,  w8_L2_N5_18= 30'h000188a1,  w8_L2_N5_19= 30'h3ff17aac,  w8_L2_N5_20= 30'h000527eb,  w8_L2_N5_21= 30'h000922f2,  w8_L2_N5_22= 30'h00000000,  w8_L2_N5_23= 30'h00000000,  w8_L2_N5_24= 30'h0009c2d7,  w8_L2_N5_25= 30'h3fff27e4,  w8_L2_N5_26= 30'h000db4e1,  w8_L2_N5_27= 30'h3ffdb960,  w8_L2_N5_28= 30'h0003a7e6,  w8_L2_N5_29= 30'h3ff69221;
reg [29:0] w8_L2_N5_30= 30'h00000000,  w8_L2_N5_31= 30'h00036ead,  w8_L2_N5_32= 30'h00091b0e,  w8_L2_N5_33= 30'h00000000,  w8_L2_N5_34= 30'h0000c106,  w8_L2_N5_35= 30'h3fffa363,  w8_L2_N5_36= 30'h00000000,  w8_L2_N5_37= 30'h00000000,  w8_L2_N5_38= 30'h3fffb636,  w8_L2_N5_39= 30'h000842bb,  w8_L2_N5_40= 30'h00037032,  w8_L2_N5_41= 30'h0000fe49,  w8_L2_N5_42= 30'h000176a0,  w8_L2_N5_43= 30'h00011f49,  w8_L2_N5_44= 30'h3ff29464,  w8_L2_N5_45= 30'h00022ea5,  w8_L2_N5_46= 30'h00041f83,  w8_L2_N5_47= 30'h3ffddda0,  w8_L2_N5_48= 30'h00000000,  w8_L2_N5_49= 30'h0009729f,  w8_L2_N5_50= 30'h00000000,  w8_L2_N5_51= 30'h3feed5d1,  w8_L2_N5_52= 30'h3ffe62fd,  w8_L2_N5_53= 30'h3ffd7d9f,  w8_L2_N5_54= 30'h00025bd7,  w8_L2_N5_55= 30'h000bdb43,  w8_L2_N5_56= 30'h00000000,  w8_L2_N5_57= 30'h00083cdd,  w8_L2_N5_58= 30'h00104ca2,  w8_L2_N5_59= 30'h0000a25f;
reg [29:0] w8_L2_N6_0= 30'h00000000,  w8_L2_N6_1= 30'h00000000,  w8_L2_N6_2= 30'h00000000,  w8_L2_N6_3= 30'h00000000,  w8_L2_N6_4= 30'h00000000,  w8_L2_N6_5= 30'h00000000,  w8_L2_N6_6= 30'h00000000,  w8_L2_N6_7= 30'h00000000,  w8_L2_N6_8= 30'h00000000,  w8_L2_N6_9= 30'h00000000,  w8_L2_N6_10= 30'h00000000,  w8_L2_N6_11= 30'h00000000,  w8_L2_N6_12= 30'h00000000,  w8_L2_N6_13= 30'h00000000,  w8_L2_N6_14= 30'h00000000,  w8_L2_N6_15= 30'h00000000,  w8_L2_N6_16= 30'h00000000,  w8_L2_N6_17= 30'h00000000,  w8_L2_N6_18= 30'h00000000,  w8_L2_N6_19= 30'h00000000,  w8_L2_N6_20= 30'h00000000,  w8_L2_N6_21= 30'h00000000,  w8_L2_N6_22= 30'h00000000,  w8_L2_N6_23= 30'h00000000,  w8_L2_N6_24= 30'h00000000,  w8_L2_N6_25= 30'h00000000,  w8_L2_N6_26= 30'h00000000,  w8_L2_N6_27= 30'h00000000,  w8_L2_N6_28= 30'h00000000,  w8_L2_N6_29= 30'h00000000;
reg [29:0] w8_L2_N6_30= 30'h00000000,  w8_L2_N6_31= 30'h00000000,  w8_L2_N6_32= 30'h00000000,  w8_L2_N6_33= 30'h00000000,  w8_L2_N6_34= 30'h00000000,  w8_L2_N6_35= 30'h00000000,  w8_L2_N6_36= 30'h00000000,  w8_L2_N6_37= 30'h00000000,  w8_L2_N6_38= 30'h00000000,  w8_L2_N6_39= 30'h00000000,  w8_L2_N6_40= 30'h00000000,  w8_L2_N6_41= 30'h00000000,  w8_L2_N6_42= 30'h00000000,  w8_L2_N6_43= 30'h00000000,  w8_L2_N6_44= 30'h00000000,  w8_L2_N6_45= 30'h00000000,  w8_L2_N6_46= 30'h00000000,  w8_L2_N6_47= 30'h00000000,  w8_L2_N6_48= 30'h00000000,  w8_L2_N6_49= 30'h00000000,  w8_L2_N6_50= 30'h00000000,  w8_L2_N6_51= 30'h00000000,  w8_L2_N6_52= 30'h00000000,  w8_L2_N6_53= 30'h00000000,  w8_L2_N6_54= 30'h00000000,  w8_L2_N6_55= 30'h00000000,  w8_L2_N6_56= 30'h00000000,  w8_L2_N6_57= 30'h00000000,  w8_L2_N6_58= 30'h00000000,  w8_L2_N6_59= 30'h00000000;
reg [29:0] w8_L2_N7_0= 30'h00000000,  w8_L2_N7_1= 30'h00000000,  w8_L2_N7_2= 30'h3ffe9b78,  w8_L2_N7_3= 30'h3ffba1a6,  w8_L2_N7_4= 30'h00000000,  w8_L2_N7_5= 30'h00000000,  w8_L2_N7_6= 30'h00000000,  w8_L2_N7_7= 30'h0007eaf0,  w8_L2_N7_8= 30'h3ff9b582,  w8_L2_N7_9= 30'h00046e79,  w8_L2_N7_10= 30'h00091ddc,  w8_L2_N7_11= 30'h00000000,  w8_L2_N7_12= 30'h3ffd8d56,  w8_L2_N7_13= 30'h3ffdb8ba,  w8_L2_N7_14= 30'h3fff22fd,  w8_L2_N7_15= 30'h00000000,  w8_L2_N7_16= 30'h3fffdf23,  w8_L2_N7_17= 30'h00000000,  w8_L2_N7_18= 30'h00047235,  w8_L2_N7_19= 30'h3ff84d7d,  w8_L2_N7_20= 30'h000272db,  w8_L2_N7_21= 30'h000aa541,  w8_L2_N7_22= 30'h00000000,  w8_L2_N7_23= 30'h00000000,  w8_L2_N7_24= 30'h000835f0,  w8_L2_N7_25= 30'h3ffffbf7,  w8_L2_N7_26= 30'h000be59a,  w8_L2_N7_27= 30'h3fff3c7e,  w8_L2_N7_28= 30'h0005a078,  w8_L2_N7_29= 30'h3ff80f67;
reg [29:0] w8_L2_N7_30= 30'h00000000,  w8_L2_N7_31= 30'h0001c377,  w8_L2_N7_32= 30'h000f753f,  w8_L2_N7_33= 30'h00004cca,  w8_L2_N7_34= 30'h00001800,  w8_L2_N7_35= 30'h3fff4385,  w8_L2_N7_36= 30'h00002072,  w8_L2_N7_37= 30'h00000000,  w8_L2_N7_38= 30'h000047d9,  w8_L2_N7_39= 30'h0009569f,  w8_L2_N7_40= 30'h0002316f,  w8_L2_N7_41= 30'h3fff1ea1,  w8_L2_N7_42= 30'h00012591,  w8_L2_N7_43= 30'h3fff5d4c,  w8_L2_N7_44= 30'h3ff67048,  w8_L2_N7_45= 30'h0003fb7c,  w8_L2_N7_46= 30'h00018767,  w8_L2_N7_47= 30'h0001b3ff,  w8_L2_N7_48= 30'h00000000,  w8_L2_N7_49= 30'h0008243f,  w8_L2_N7_50= 30'h00000000,  w8_L2_N7_51= 30'h3ff8352b,  w8_L2_N7_52= 30'h00035baa,  w8_L2_N7_53= 30'h3fff81b0,  w8_L2_N7_54= 30'h000208ee,  w8_L2_N7_55= 30'h000d56c4,  w8_L2_N7_56= 30'h3ffff75a,  w8_L2_N7_57= 30'h00068b0d,  w8_L2_N7_58= 30'h000d4e96,  w8_L2_N7_59= 30'h00045b79;
reg [29:0] w8_L2_N8_0= 30'h00000000,  w8_L2_N8_1= 30'h00000000,  w8_L2_N8_2= 30'h00000000,  w8_L2_N8_3= 30'h00000000,  w8_L2_N8_4= 30'h00000000,  w8_L2_N8_5= 30'h00000000,  w8_L2_N8_6= 30'h00000000,  w8_L2_N8_7= 30'h00000000,  w8_L2_N8_8= 30'h00000000,  w8_L2_N8_9= 30'h00000000,  w8_L2_N8_10= 30'h00000000,  w8_L2_N8_11= 30'h00000000,  w8_L2_N8_12= 30'h00000000,  w8_L2_N8_13= 30'h00000000,  w8_L2_N8_14= 30'h00000000,  w8_L2_N8_15= 30'h00000000,  w8_L2_N8_16= 30'h00000000,  w8_L2_N8_17= 30'h00000000,  w8_L2_N8_18= 30'h00000000,  w8_L2_N8_19= 30'h00000000,  w8_L2_N8_20= 30'h00000000,  w8_L2_N8_21= 30'h00000000,  w8_L2_N8_22= 30'h00000000,  w8_L2_N8_23= 30'h00000000,  w8_L2_N8_24= 30'h00000000,  w8_L2_N8_25= 30'h00000000,  w8_L2_N8_26= 30'h00000000,  w8_L2_N8_27= 30'h00000000,  w8_L2_N8_28= 30'h00000000,  w8_L2_N8_29= 30'h00000000;
reg [29:0] w8_L2_N8_30= 30'h00000000,  w8_L2_N8_31= 30'h00000000,  w8_L2_N8_32= 30'h00000000,  w8_L2_N8_33= 30'h00000000,  w8_L2_N8_34= 30'h00000000,  w8_L2_N8_35= 30'h00000000,  w8_L2_N8_36= 30'h00000000,  w8_L2_N8_37= 30'h00000000,  w8_L2_N8_38= 30'h00000000,  w8_L2_N8_39= 30'h00000000,  w8_L2_N8_40= 30'h00000000,  w8_L2_N8_41= 30'h00000000,  w8_L2_N8_42= 30'h00000000,  w8_L2_N8_43= 30'h00000000,  w8_L2_N8_44= 30'h00000000,  w8_L2_N8_45= 30'h00000000,  w8_L2_N8_46= 30'h00000000,  w8_L2_N8_47= 30'h00000000,  w8_L2_N8_48= 30'h00000000,  w8_L2_N8_49= 30'h00000000,  w8_L2_N8_50= 30'h00000000,  w8_L2_N8_51= 30'h00000000,  w8_L2_N8_52= 30'h00000000,  w8_L2_N8_53= 30'h00000000,  w8_L2_N8_54= 30'h00000000,  w8_L2_N8_55= 30'h00000000,  w8_L2_N8_56= 30'h00000000,  w8_L2_N8_57= 30'h00000000,  w8_L2_N8_58= 30'h00000000,  w8_L2_N8_59= 30'h00000000;
reg [29:0] w8_L2_N9_0= 30'h00000000,  w8_L2_N9_1= 30'h00000000,  w8_L2_N9_2= 30'h000136a6,  w8_L2_N9_3= 30'h000430d3,  w8_L2_N9_4= 30'h00000000,  w8_L2_N9_5= 30'h00000000,  w8_L2_N9_6= 30'h00000000,  w8_L2_N9_7= 30'h3ffecc99,  w8_L2_N9_8= 30'h3ffeddfd,  w8_L2_N9_9= 30'h00014873,  w8_L2_N9_10= 30'h3fff34df,  w8_L2_N9_11= 30'h00000000,  w8_L2_N9_12= 30'h00020916,  w8_L2_N9_13= 30'h3fffb0f0,  w8_L2_N9_14= 30'h000280b6,  w8_L2_N9_15= 30'h00000000,  w8_L2_N9_16= 30'h3ffffff9,  w8_L2_N9_17= 30'h00000000,  w8_L2_N9_18= 30'h00012a8c,  w8_L2_N9_19= 30'h3fff0cd0,  w8_L2_N9_20= 30'h3fff539e,  w8_L2_N9_21= 30'h3ffdb64b,  w8_L2_N9_22= 30'h00000000,  w8_L2_N9_23= 30'h00000000,  w8_L2_N9_24= 30'h0000102c,  w8_L2_N9_25= 30'h3ffffa39,  w8_L2_N9_26= 30'h3ffebff8,  w8_L2_N9_27= 30'h00035956,  w8_L2_N9_28= 30'h3fff1994,  w8_L2_N9_29= 30'h0001279b;
reg [29:0] w8_L2_N9_30= 30'h00000000,  w8_L2_N9_31= 30'h0002c15e,  w8_L2_N9_32= 30'h3ffe351b,  w8_L2_N9_33= 30'h3ffff054,  w8_L2_N9_34= 30'h00032d84,  w8_L2_N9_35= 30'h0002f679,  w8_L2_N9_36= 30'h3fffffe0,  w8_L2_N9_37= 30'h00000000,  w8_L2_N9_38= 30'h0003f98a,  w8_L2_N9_39= 30'h3fffac52,  w8_L2_N9_40= 30'h00017d57,  w8_L2_N9_41= 30'h000203db,  w8_L2_N9_42= 30'h0000a527,  w8_L2_N9_43= 30'h0002db1d,  w8_L2_N9_44= 30'h3fff7f93,  w8_L2_N9_45= 30'h0000a348,  w8_L2_N9_46= 30'h00006ed3,  w8_L2_N9_47= 30'h0000ae22,  w8_L2_N9_48= 30'h00000000,  w8_L2_N9_49= 30'h3ffd62ad,  w8_L2_N9_50= 30'h00000000,  w8_L2_N9_51= 30'h3fff7056,  w8_L2_N9_52= 30'h3ffe1f51,  w8_L2_N9_53= 30'h00030412,  w8_L2_N9_54= 30'h00017157,  w8_L2_N9_55= 30'h3ffdebf4,  w8_L2_N9_56= 30'h00000005,  w8_L2_N9_57= 30'h00004f70,  w8_L2_N9_58= 30'h3ffed48c,  w8_L2_N9_59= 30'h0002945e;
reg [29:0] w8_L2_N10_0= 30'h00000000,  w8_L2_N10_1= 30'h00000000,  w8_L2_N10_2= 30'h00000000,  w8_L2_N10_3= 30'h00000000,  w8_L2_N10_4= 30'h00000000,  w8_L2_N10_5= 30'h00000000,  w8_L2_N10_6= 30'h00000000,  w8_L2_N10_7= 30'h00000000,  w8_L2_N10_8= 30'h00000000,  w8_L2_N10_9= 30'h00000000,  w8_L2_N10_10= 30'h00000000,  w8_L2_N10_11= 30'h00000000,  w8_L2_N10_12= 30'h00000000,  w8_L2_N10_13= 30'h00000000,  w8_L2_N10_14= 30'h00000000,  w8_L2_N10_15= 30'h00000000,  w8_L2_N10_16= 30'h00000000,  w8_L2_N10_17= 30'h00000000,  w8_L2_N10_18= 30'h00000000,  w8_L2_N10_19= 30'h00000000,  w8_L2_N10_20= 30'h00000000,  w8_L2_N10_21= 30'h00000000,  w8_L2_N10_22= 30'h00000000,  w8_L2_N10_23= 30'h00000000,  w8_L2_N10_24= 30'h00000000,  w8_L2_N10_25= 30'h00000000,  w8_L2_N10_26= 30'h00000000,  w8_L2_N10_27= 30'h00000000,  w8_L2_N10_28= 30'h00000000,  w8_L2_N10_29= 30'h00000000;
reg [29:0] w8_L2_N10_30= 30'h00000000,  w8_L2_N10_31= 30'h00000000,  w8_L2_N10_32= 30'h00000000,  w8_L2_N10_33= 30'h00000000,  w8_L2_N10_34= 30'h00000000,  w8_L2_N10_35= 30'h00000000,  w8_L2_N10_36= 30'h00000000,  w8_L2_N10_37= 30'h00000000,  w8_L2_N10_38= 30'h00000000,  w8_L2_N10_39= 30'h00000000,  w8_L2_N10_40= 30'h00000000,  w8_L2_N10_41= 30'h00000000,  w8_L2_N10_42= 30'h00000000,  w8_L2_N10_43= 30'h00000000,  w8_L2_N10_44= 30'h00000000,  w8_L2_N10_45= 30'h00000000,  w8_L2_N10_46= 30'h00000000,  w8_L2_N10_47= 30'h00000000,  w8_L2_N10_48= 30'h00000000,  w8_L2_N10_49= 30'h00000000,  w8_L2_N10_50= 30'h00000000,  w8_L2_N10_51= 30'h00000000,  w8_L2_N10_52= 30'h00000000,  w8_L2_N10_53= 30'h00000000,  w8_L2_N10_54= 30'h00000000,  w8_L2_N10_55= 30'h00000000,  w8_L2_N10_56= 30'h00000000,  w8_L2_N10_57= 30'h00000000,  w8_L2_N10_58= 30'h00000000,  w8_L2_N10_59= 30'h00000000;
reg [29:0] w8_L2_N11_0= 30'h00000000,  w8_L2_N11_1= 30'h00000000,  w8_L2_N11_2= 30'h3ffeea38,  w8_L2_N11_3= 30'h00000000,  w8_L2_N11_4= 30'h00000000,  w8_L2_N11_5= 30'h00000000,  w8_L2_N11_6= 30'h00000000,  w8_L2_N11_7= 30'h0000c210,  w8_L2_N11_8= 30'h00000f86,  w8_L2_N11_9= 30'h00001126,  w8_L2_N11_10= 30'h00000f43,  w8_L2_N11_11= 30'h00000000,  w8_L2_N11_12= 30'h00000000,  w8_L2_N11_13= 30'h00000000,  w8_L2_N11_14= 30'h0000c108,  w8_L2_N11_15= 30'h00000000,  w8_L2_N11_16= 30'h3fff4eb1,  w8_L2_N11_17= 30'h00000000,  w8_L2_N11_18= 30'h000056e0,  w8_L2_N11_19= 30'h3fff50fb,  w8_L2_N11_20= 30'h00001dba,  w8_L2_N11_21= 30'h00009b1f,  w8_L2_N11_22= 30'h00000000,  w8_L2_N11_23= 30'h00000000,  w8_L2_N11_24= 30'h00000000,  w8_L2_N11_25= 30'h0000d2d5,  w8_L2_N11_26= 30'h3ffe96ca,  w8_L2_N11_27= 30'h3ffee06d,  w8_L2_N11_28= 30'h0000d846,  w8_L2_N11_29= 30'h3fff1120;
reg [29:0] w8_L2_N11_30= 30'h00000000,  w8_L2_N11_31= 30'h00000000,  w8_L2_N11_32= 30'h3ffffe78,  w8_L2_N11_33= 30'h00003897,  w8_L2_N11_34= 30'h00000000,  w8_L2_N11_35= 30'h3fffe111,  w8_L2_N11_36= 30'h3fffd67f,  w8_L2_N11_37= 30'h00000000,  w8_L2_N11_38= 30'h00008595,  w8_L2_N11_39= 30'h3fffbbae,  w8_L2_N11_40= 30'h3ffe555c,  w8_L2_N11_41= 30'h00000000,  w8_L2_N11_42= 30'h3fff95cc,  w8_L2_N11_43= 30'h00000468,  w8_L2_N11_44= 30'h3fff727c,  w8_L2_N11_45= 30'h000001d7,  w8_L2_N11_46= 30'h00004862,  w8_L2_N11_47= 30'h000004ff,  w8_L2_N11_48= 30'h3ffffff8,  w8_L2_N11_49= 30'h3fff3b89,  w8_L2_N11_50= 30'h00000000,  w8_L2_N11_51= 30'h00000028,  w8_L2_N11_52= 30'h00000000,  w8_L2_N11_53= 30'h3fffa0e5,  w8_L2_N11_54= 30'h00005029,  w8_L2_N11_55= 30'h3fffdb5d,  w8_L2_N11_56= 30'h3fff9599,  w8_L2_N11_57= 30'h00000000,  w8_L2_N11_58= 30'h0000e3ee,  w8_L2_N11_59= 30'h00000fc5;
reg [29:0] w8_L2_N12_0= 30'h00000000,  w8_L2_N12_1= 30'h00000000,  w8_L2_N12_2= 30'h3fffb9a0,  w8_L2_N12_3= 30'h3fffcd95,  w8_L2_N12_4= 30'h00000000,  w8_L2_N12_5= 30'h00000000,  w8_L2_N12_6= 30'h00000000,  w8_L2_N12_7= 30'h3fffffc0,  w8_L2_N12_8= 30'h0000081c,  w8_L2_N12_9= 30'h3fffdc35,  w8_L2_N12_10= 30'h00000049,  w8_L2_N12_11= 30'h00000000,  w8_L2_N12_12= 30'h3fffb7f7,  w8_L2_N12_13= 30'h00000001,  w8_L2_N12_14= 30'h3fffc47a,  w8_L2_N12_15= 30'h00000000,  w8_L2_N12_16= 30'h00000000,  w8_L2_N12_17= 30'h00000000,  w8_L2_N12_18= 30'h3fffe878,  w8_L2_N12_19= 30'h00000379,  w8_L2_N12_20= 30'h3fffe7cb,  w8_L2_N12_21= 30'h3ffffec5,  w8_L2_N12_22= 30'h00000000,  w8_L2_N12_23= 30'h00000000,  w8_L2_N12_24= 30'h3ffffa07,  w8_L2_N12_25= 30'h3fffee8b,  w8_L2_N12_26= 30'h00000004,  w8_L2_N12_27= 30'h3fffa3ee,  w8_L2_N12_28= 30'h00000065,  w8_L2_N12_29= 30'h3fffffb8;
reg [29:0] w8_L2_N12_30= 30'h00000000,  w8_L2_N12_31= 30'h3fffc1d3,  w8_L2_N12_32= 30'h00000005,  w8_L2_N12_33= 30'h00000000,  w8_L2_N12_34= 30'h3fffc25c,  w8_L2_N12_35= 30'h3fffc418,  w8_L2_N12_36= 30'h00000000,  w8_L2_N12_37= 30'h00000000,  w8_L2_N12_38= 30'h3fffc83c,  w8_L2_N12_39= 30'h3ffffa40,  w8_L2_N12_40= 30'h3fffb7f1,  w8_L2_N12_41= 30'h3fffc07b,  w8_L2_N12_42= 30'h3fffd65a,  w8_L2_N12_43= 30'h3fffbf84,  w8_L2_N12_44= 30'h0000019c,  w8_L2_N12_45= 30'h3fffd613,  w8_L2_N12_46= 30'h3ffff8b8,  w8_L2_N12_47= 30'h3fffdde9,  w8_L2_N12_48= 30'h00000000,  w8_L2_N12_49= 30'h00000205,  w8_L2_N12_50= 30'h00000000,  w8_L2_N12_51= 30'h00000568,  w8_L2_N12_52= 30'h0000022f,  w8_L2_N12_53= 30'h3fffb9f9,  w8_L2_N12_54= 30'h3fffc2c5,  w8_L2_N12_55= 30'h3fffffde,  w8_L2_N12_56= 30'h00000000,  w8_L2_N12_57= 30'h3ffff070,  w8_L2_N12_58= 30'h00000001,  w8_L2_N12_59= 30'h3fffd843;
reg [29:0] w8_L2_N13_0= 30'h00000000,  w8_L2_N13_1= 30'h00000000,  w8_L2_N13_2= 30'h00000000,  w8_L2_N13_3= 30'h00000000,  w8_L2_N13_4= 30'h00000000,  w8_L2_N13_5= 30'h00000000,  w8_L2_N13_6= 30'h00000000,  w8_L2_N13_7= 30'h00000000,  w8_L2_N13_8= 30'h00000000,  w8_L2_N13_9= 30'h00000000,  w8_L2_N13_10= 30'h00000000,  w8_L2_N13_11= 30'h00000000,  w8_L2_N13_12= 30'h00000000,  w8_L2_N13_13= 30'h00000000,  w8_L2_N13_14= 30'h00000000,  w8_L2_N13_15= 30'h00000000,  w8_L2_N13_16= 30'h00000000,  w8_L2_N13_17= 30'h00000000,  w8_L2_N13_18= 30'h00000000,  w8_L2_N13_19= 30'h00000000,  w8_L2_N13_20= 30'h00000000,  w8_L2_N13_21= 30'h00000000,  w8_L2_N13_22= 30'h00000000,  w8_L2_N13_23= 30'h00000000,  w8_L2_N13_24= 30'h00000000,  w8_L2_N13_25= 30'h00000000,  w8_L2_N13_26= 30'h00000000,  w8_L2_N13_27= 30'h00000000,  w8_L2_N13_28= 30'h00000000,  w8_L2_N13_29= 30'h00000000;
reg [29:0] w8_L2_N13_30= 30'h00000000,  w8_L2_N13_31= 30'h00000000,  w8_L2_N13_32= 30'h00000000,  w8_L2_N13_33= 30'h00000000,  w8_L2_N13_34= 30'h00000000,  w8_L2_N13_35= 30'h00000000,  w8_L2_N13_36= 30'h00000000,  w8_L2_N13_37= 30'h00000000,  w8_L2_N13_38= 30'h00000000,  w8_L2_N13_39= 30'h00000000,  w8_L2_N13_40= 30'h00000000,  w8_L2_N13_41= 30'h00000000,  w8_L2_N13_42= 30'h00000000,  w8_L2_N13_43= 30'h00000000,  w8_L2_N13_44= 30'h00000000,  w8_L2_N13_45= 30'h00000000,  w8_L2_N13_46= 30'h00000000,  w8_L2_N13_47= 30'h00000000,  w8_L2_N13_48= 30'h00000000,  w8_L2_N13_49= 30'h00000000,  w8_L2_N13_50= 30'h00000000,  w8_L2_N13_51= 30'h00000000,  w8_L2_N13_52= 30'h00000000,  w8_L2_N13_53= 30'h00000000,  w8_L2_N13_54= 30'h00000000,  w8_L2_N13_55= 30'h00000000,  w8_L2_N13_56= 30'h00000000,  w8_L2_N13_57= 30'h00000000,  w8_L2_N13_58= 30'h00000000,  w8_L2_N13_59= 30'h00000000;
reg [29:0] w8_L2_N14_0= 30'h00000000,  w8_L2_N14_1= 30'h00000000,  w8_L2_N14_2= 30'h00000000,  w8_L2_N14_3= 30'h00000000,  w8_L2_N14_4= 30'h00000000,  w8_L2_N14_5= 30'h00000000,  w8_L2_N14_6= 30'h00000000,  w8_L2_N14_7= 30'h00000000,  w8_L2_N14_8= 30'h00000000,  w8_L2_N14_9= 30'h00000000,  w8_L2_N14_10= 30'h00000000,  w8_L2_N14_11= 30'h00000000,  w8_L2_N14_12= 30'h00000000,  w8_L2_N14_13= 30'h00000000,  w8_L2_N14_14= 30'h00000000,  w8_L2_N14_15= 30'h00000000,  w8_L2_N14_16= 30'h00000000,  w8_L2_N14_17= 30'h00000000,  w8_L2_N14_18= 30'h00000000,  w8_L2_N14_19= 30'h00000000,  w8_L2_N14_20= 30'h00000000,  w8_L2_N14_21= 30'h00000000,  w8_L2_N14_22= 30'h00000000,  w8_L2_N14_23= 30'h00000000,  w8_L2_N14_24= 30'h00000000,  w8_L2_N14_25= 30'h00000000,  w8_L2_N14_26= 30'h00000000,  w8_L2_N14_27= 30'h00000000,  w8_L2_N14_28= 30'h00000000,  w8_L2_N14_29= 30'h00000000;
reg [29:0] w8_L2_N14_30= 30'h00000000,  w8_L2_N14_31= 30'h00000000,  w8_L2_N14_32= 30'h00000000,  w8_L2_N14_33= 30'h00000000,  w8_L2_N14_34= 30'h00000000,  w8_L2_N14_35= 30'h00000000,  w8_L2_N14_36= 30'h00000000,  w8_L2_N14_37= 30'h00000000,  w8_L2_N14_38= 30'h00000000,  w8_L2_N14_39= 30'h00000000,  w8_L2_N14_40= 30'h00000000,  w8_L2_N14_41= 30'h00000000,  w8_L2_N14_42= 30'h00000000,  w8_L2_N14_43= 30'h00000000,  w8_L2_N14_44= 30'h00000000,  w8_L2_N14_45= 30'h00000000,  w8_L2_N14_46= 30'h00000000,  w8_L2_N14_47= 30'h00000000,  w8_L2_N14_48= 30'h00000000,  w8_L2_N14_49= 30'h00000000,  w8_L2_N14_50= 30'h00000000,  w8_L2_N14_51= 30'h00000000,  w8_L2_N14_52= 30'h00000000,  w8_L2_N14_53= 30'h00000000,  w8_L2_N14_54= 30'h00000000,  w8_L2_N14_55= 30'h00000000,  w8_L2_N14_56= 30'h00000000,  w8_L2_N14_57= 30'h00000000,  w8_L2_N14_58= 30'h00000000,  w8_L2_N14_59= 30'h00000000;
reg [29:0] w8_L2_N15_0= 30'h00000000,  w8_L2_N15_1= 30'h00000000,  w8_L2_N15_2= 30'h3ffc9f08,  w8_L2_N15_3= 30'h3ffc88ef,  w8_L2_N15_4= 30'h00000000,  w8_L2_N15_5= 30'h00000000,  w8_L2_N15_6= 30'h00000000,  w8_L2_N15_7= 30'h00040dd3,  w8_L2_N15_8= 30'h3fff52be,  w8_L2_N15_9= 30'h0002f15e,  w8_L2_N15_10= 30'h000586b5,  w8_L2_N15_11= 30'h00000000,  w8_L2_N15_12= 30'h3ffcdd1e,  w8_L2_N15_13= 30'h0001712d,  w8_L2_N15_14= 30'h00026dde,  w8_L2_N15_15= 30'h00000000,  w8_L2_N15_16= 30'h3fff5df4,  w8_L2_N15_17= 30'h00000000,  w8_L2_N15_18= 30'h000061b6,  w8_L2_N15_19= 30'h3fff03ce,  w8_L2_N15_20= 30'h000559e0,  w8_L2_N15_21= 30'h00080e7b,  w8_L2_N15_22= 30'h00000000,  w8_L2_N15_23= 30'h00000000,  w8_L2_N15_24= 30'h000a4c28,  w8_L2_N15_25= 30'h000340f2,  w8_L2_N15_26= 30'h00069c05,  w8_L2_N15_27= 30'h00024fc4,  w8_L2_N15_28= 30'h00064a95,  w8_L2_N15_29= 30'h3ffdc429;
reg [29:0] w8_L2_N15_30= 30'h00000000,  w8_L2_N15_31= 30'h3ffd760b,  w8_L2_N15_32= 30'h000d01d1,  w8_L2_N15_33= 30'h3fff024e,  w8_L2_N15_34= 30'h3ffb3421,  w8_L2_N15_35= 30'h3ffd7007,  w8_L2_N15_36= 30'h3fffa778,  w8_L2_N15_37= 30'h00000000,  w8_L2_N15_38= 30'h3ffd4377,  w8_L2_N15_39= 30'h0005dc86,  w8_L2_N15_40= 30'h3fff3e4f,  w8_L2_N15_41= 30'h3ffddb9e,  w8_L2_N15_42= 30'h00046201,  w8_L2_N15_43= 30'h3ffc8c03,  w8_L2_N15_44= 30'h3ffe3d37,  w8_L2_N15_45= 30'h0001d59b,  w8_L2_N15_46= 30'h0004f88a,  w8_L2_N15_47= 30'h00032322,  w8_L2_N15_48= 30'h3ffffffd,  w8_L2_N15_49= 30'h00083b95,  w8_L2_N15_50= 30'h00000000,  w8_L2_N15_51= 30'h3ffc22a5,  w8_L2_N15_52= 30'h00093000,  w8_L2_N15_53= 30'h0000fda7,  w8_L2_N15_54= 30'h0001151b,  w8_L2_N15_55= 30'h000b968d,  w8_L2_N15_56= 30'h3fffcb10,  w8_L2_N15_57= 30'h00080ca4,  w8_L2_N15_58= 30'h000baf46,  w8_L2_N15_59= 30'h0001872b;
reg [29:0] w8_L2_N16_0= 30'h00000000,  w8_L2_N16_1= 30'h00000000,  w8_L2_N16_2= 30'h00000000,  w8_L2_N16_3= 30'h00000000,  w8_L2_N16_4= 30'h00000000,  w8_L2_N16_5= 30'h00000000,  w8_L2_N16_6= 30'h00000000,  w8_L2_N16_7= 30'h00000000,  w8_L2_N16_8= 30'h00000000,  w8_L2_N16_9= 30'h00000000,  w8_L2_N16_10= 30'h00000000,  w8_L2_N16_11= 30'h00000000,  w8_L2_N16_12= 30'h00000000,  w8_L2_N16_13= 30'h00000000,  w8_L2_N16_14= 30'h00000000,  w8_L2_N16_15= 30'h00000000,  w8_L2_N16_16= 30'h00000000,  w8_L2_N16_17= 30'h00000000,  w8_L2_N16_18= 30'h00000000,  w8_L2_N16_19= 30'h00000000,  w8_L2_N16_20= 30'h00000000,  w8_L2_N16_21= 30'h00000000,  w8_L2_N16_22= 30'h00000000,  w8_L2_N16_23= 30'h00000000,  w8_L2_N16_24= 30'h00000000,  w8_L2_N16_25= 30'h00000000,  w8_L2_N16_26= 30'h00000000,  w8_L2_N16_27= 30'h00000000,  w8_L2_N16_28= 30'h00000000,  w8_L2_N16_29= 30'h00000000;
reg [29:0] w8_L2_N16_30= 30'h00000000,  w8_L2_N16_31= 30'h00000000,  w8_L2_N16_32= 30'h00000000,  w8_L2_N16_33= 30'h00000000,  w8_L2_N16_34= 30'h00000000,  w8_L2_N16_35= 30'h00000000,  w8_L2_N16_36= 30'h00000000,  w8_L2_N16_37= 30'h00000000,  w8_L2_N16_38= 30'h00000000,  w8_L2_N16_39= 30'h00000000,  w8_L2_N16_40= 30'h00000000,  w8_L2_N16_41= 30'h00000000,  w8_L2_N16_42= 30'h00000000,  w8_L2_N16_43= 30'h00000000,  w8_L2_N16_44= 30'h00000000,  w8_L2_N16_45= 30'h00000000,  w8_L2_N16_46= 30'h00000000,  w8_L2_N16_47= 30'h00000000,  w8_L2_N16_48= 30'h00000000,  w8_L2_N16_49= 30'h00000000,  w8_L2_N16_50= 30'h00000000,  w8_L2_N16_51= 30'h00000000,  w8_L2_N16_52= 30'h00000000,  w8_L2_N16_53= 30'h00000000,  w8_L2_N16_54= 30'h00000000,  w8_L2_N16_55= 30'h00000000,  w8_L2_N16_56= 30'h00000000,  w8_L2_N16_57= 30'h00000000,  w8_L2_N16_58= 30'h00000000,  w8_L2_N16_59= 30'h00000000;
reg [29:0] w8_L2_N17_0= 30'h00000000,  w8_L2_N17_1= 30'h00000000,  w8_L2_N17_2= 30'h00007e81,  w8_L2_N17_3= 30'h00035848,  w8_L2_N17_4= 30'h00000000,  w8_L2_N17_5= 30'h00000000,  w8_L2_N17_6= 30'h00000000,  w8_L2_N17_7= 30'h3ffbe6b7,  w8_L2_N17_8= 30'h0001e1f0,  w8_L2_N17_9= 30'h3ffe01eb,  w8_L2_N17_10= 30'h3ffb9a94,  w8_L2_N17_11= 30'h00000000,  w8_L2_N17_12= 30'h00025bdb,  w8_L2_N17_13= 30'h00011681,  w8_L2_N17_14= 30'h00016b07,  w8_L2_N17_15= 30'h00000000,  w8_L2_N17_16= 30'h00000345,  w8_L2_N17_17= 30'h00000000,  w8_L2_N17_18= 30'h3ffe9fbf,  w8_L2_N17_19= 30'h0002b3f6,  w8_L2_N17_20= 30'h3fff7789,  w8_L2_N17_21= 30'h3ffa73c5,  w8_L2_N17_22= 30'h00000000,  w8_L2_N17_23= 30'h00000000,  w8_L2_N17_24= 30'h3ff96f74,  w8_L2_N17_25= 30'h000146ba,  w8_L2_N17_26= 30'h3ffaf49a,  w8_L2_N17_27= 30'h0002acfc,  w8_L2_N17_28= 30'h3fff65e1,  w8_L2_N17_29= 30'h0002fd6e;
reg [29:0] w8_L2_N17_30= 30'h00000000,  w8_L2_N17_31= 30'h000380f2,  w8_L2_N17_32= 30'h3ff870f5,  w8_L2_N17_33= 30'h3fff10da,  w8_L2_N17_34= 30'h00035bf1,  w8_L2_N17_35= 30'h00039a92,  w8_L2_N17_36= 30'h3fffb637,  w8_L2_N17_37= 30'h00000000,  w8_L2_N17_38= 30'h000279f5,  w8_L2_N17_39= 30'h3ff9cf38,  w8_L2_N17_40= 30'h3fffe81b,  w8_L2_N17_41= 30'h0002aeca,  w8_L2_N17_42= 30'h0001d5ce,  w8_L2_N17_43= 30'h0002b561,  w8_L2_N17_44= 30'h00053900,  w8_L2_N17_45= 30'h00004cca,  w8_L2_N17_46= 30'h00007e8c,  w8_L2_N17_47= 30'h0001c444,  w8_L2_N17_48= 30'h00000002,  w8_L2_N17_49= 30'h3ffa210e,  w8_L2_N17_50= 30'h00000000,  w8_L2_N17_51= 30'h00026713,  w8_L2_N17_52= 30'h3ffb10a6,  w8_L2_N17_53= 30'h0000946f,  w8_L2_N17_54= 30'h000281da,  w8_L2_N17_55= 30'h3ff94283,  w8_L2_N17_56= 30'h000039ed,  w8_L2_N17_57= 30'h3ffb560b,  w8_L2_N17_58= 30'h3ffa960b,  w8_L2_N17_59= 30'h3ffd8ef4;
reg [29:0] w8_L2_N18_0= 30'h00000000,  w8_L2_N18_1= 30'h00000000,  w8_L2_N18_2= 30'h3ffe50d0,  w8_L2_N18_3= 30'h3ffdf035,  w8_L2_N18_4= 30'h00000000,  w8_L2_N18_5= 30'h00000000,  w8_L2_N18_6= 30'h00000000,  w8_L2_N18_7= 30'h000399f3,  w8_L2_N18_8= 30'h000420f7,  w8_L2_N18_9= 30'h0001c02b,  w8_L2_N18_10= 30'h000465e0,  w8_L2_N18_11= 30'h00000000,  w8_L2_N18_12= 30'h3ffa6b7a,  w8_L2_N18_13= 30'h000532b3,  w8_L2_N18_14= 30'h3fff3fb0,  w8_L2_N18_15= 30'h00000000,  w8_L2_N18_16= 30'h00000dee,  w8_L2_N18_17= 30'h00000000,  w8_L2_N18_18= 30'h0000b37a,  w8_L2_N18_19= 30'h00043d79,  w8_L2_N18_20= 30'h0001455a,  w8_L2_N18_21= 30'h00055cb2,  w8_L2_N18_22= 30'h00000000,  w8_L2_N18_23= 30'h00000000,  w8_L2_N18_24= 30'h0000a432,  w8_L2_N18_25= 30'h00022524,  w8_L2_N18_26= 30'h00039010,  w8_L2_N18_27= 30'h3fff9451,  w8_L2_N18_28= 30'h00055341,  w8_L2_N18_29= 30'h000247fc;
reg [29:0] w8_L2_N18_30= 30'h00000000,  w8_L2_N18_31= 30'h3ffea416,  w8_L2_N18_32= 30'h00040abe,  w8_L2_N18_33= 30'h3fffefa0,  w8_L2_N18_34= 30'h3ffd50f1,  w8_L2_N18_35= 30'h3ffc5949,  w8_L2_N18_36= 30'h3fffe38b,  w8_L2_N18_37= 30'h00000000,  w8_L2_N18_38= 30'h3ffbf5e5,  w8_L2_N18_39= 30'h3ffea087,  w8_L2_N18_40= 30'h0000b620,  w8_L2_N18_41= 30'h3ffafe8d,  w8_L2_N18_42= 30'h0002bd7a,  w8_L2_N18_43= 30'h3ffc0fb6,  w8_L2_N18_44= 30'h00046749,  w8_L2_N18_45= 30'h0000c0ed,  w8_L2_N18_46= 30'h0004ce40,  w8_L2_N18_47= 30'h00003201,  w8_L2_N18_48= 30'h00000000,  w8_L2_N18_49= 30'h00033fdf,  w8_L2_N18_50= 30'h00000000,  w8_L2_N18_51= 30'h00060fda,  w8_L2_N18_52= 30'h000c68d1,  w8_L2_N18_53= 30'h3ffd4cb9,  w8_L2_N18_54= 30'h3fff2294,  w8_L2_N18_55= 30'h0004245f,  w8_L2_N18_56= 30'h0000000a,  w8_L2_N18_57= 30'h000019f6,  w8_L2_N18_58= 30'h00028425,  w8_L2_N18_59= 30'h3fff88ea;
reg [29:0] w8_L2_N19_0= 30'h00000000,  w8_L2_N19_1= 30'h00000000,  w8_L2_N19_2= 30'h00006b91,  w8_L2_N19_3= 30'h0003f5f6,  w8_L2_N19_4= 30'h00000000,  w8_L2_N19_5= 30'h00000000,  w8_L2_N19_6= 30'h00000000,  w8_L2_N19_7= 30'h3ffc2478,  w8_L2_N19_8= 30'h00061391,  w8_L2_N19_9= 30'h3ffe5a97,  w8_L2_N19_10= 30'h3ff864fe,  w8_L2_N19_11= 30'h00000000,  w8_L2_N19_12= 30'h0000aaca,  w8_L2_N19_13= 30'h00013fdb,  w8_L2_N19_14= 30'h0001e77d,  w8_L2_N19_15= 30'h00000000,  w8_L2_N19_16= 30'h0000864b,  w8_L2_N19_17= 30'h00000000,  w8_L2_N19_18= 30'h3ffed9d5,  w8_L2_N19_19= 30'h00077d44,  w8_L2_N19_20= 30'h3ffc7e6a,  w8_L2_N19_21= 30'h3ff7ed0c,  w8_L2_N19_22= 30'h00000000,  w8_L2_N19_23= 30'h00000000,  w8_L2_N19_24= 30'h3ff75478,  w8_L2_N19_25= 30'h0001d72c,  w8_L2_N19_26= 30'h3ff653a8,  w8_L2_N19_27= 30'h00008f75,  w8_L2_N19_28= 30'h3ffc6fc0,  w8_L2_N19_29= 30'h0006b532;
reg [29:0] w8_L2_N19_30= 30'h00000000,  w8_L2_N19_31= 30'h3fff6958,  w8_L2_N19_32= 30'h3ff0a863,  w8_L2_N19_33= 30'h00009dd8,  w8_L2_N19_34= 30'h0002a38d,  w8_L2_N19_35= 30'h0001d0a3,  w8_L2_N19_36= 30'h000001f1,  w8_L2_N19_37= 30'h00000000,  w8_L2_N19_38= 30'h00027571,  w8_L2_N19_39= 30'h3ffa45c4,  w8_L2_N19_40= 30'h000027bc,  w8_L2_N19_41= 30'h00013727,  w8_L2_N19_42= 30'h3ffff6ac,  w8_L2_N19_43= 30'h0001cbe8,  w8_L2_N19_44= 30'h0009cc6b,  w8_L2_N19_45= 30'h3ffcc08d,  w8_L2_N19_46= 30'h3ffc1e78,  w8_L2_N19_47= 30'h00019663,  w8_L2_N19_48= 30'h00000023,  w8_L2_N19_49= 30'h3ff5fd7e,  w8_L2_N19_50= 30'h00000000,  w8_L2_N19_51= 30'h000bf8f4,  w8_L2_N19_52= 30'h3ffa6b3e,  w8_L2_N19_53= 30'h0001b83c,  w8_L2_N19_54= 30'h000136e8,  w8_L2_N19_55= 30'h3ff1e662,  w8_L2_N19_56= 30'h000006c1,  w8_L2_N19_57= 30'h3ff67910,  w8_L2_N19_58= 30'h3ff5eafe,  w8_L2_N19_59= 30'h3ffc68db;
reg [29:0] w8_L2_N20_0= 30'h00000000,  w8_L2_N20_1= 30'h00000000,  w8_L2_N20_2= 30'h3fffd4ce,  w8_L2_N20_3= 30'h3ffd1538,  w8_L2_N20_4= 30'h00000000,  w8_L2_N20_5= 30'h00000000,  w8_L2_N20_6= 30'h00000000,  w8_L2_N20_7= 30'h00059725,  w8_L2_N20_8= 30'h3ff465fa,  w8_L2_N20_9= 30'h000253d8,  w8_L2_N20_10= 30'h00067739,  w8_L2_N20_11= 30'h00000000,  w8_L2_N20_12= 30'h0001ace1,  w8_L2_N20_13= 30'h3ffbebda,  w8_L2_N20_14= 30'h00015154,  w8_L2_N20_15= 30'h00000000,  w8_L2_N20_16= 30'h00000012,  w8_L2_N20_17= 30'h00000000,  w8_L2_N20_18= 30'h000285a9,  w8_L2_N20_19= 30'h3ff40d6e,  w8_L2_N20_20= 30'h00013263,  w8_L2_N20_21= 30'h0006543e,  w8_L2_N20_22= 30'h00000000,  w8_L2_N20_23= 30'h00000000,  w8_L2_N20_24= 30'h000894f8,  w8_L2_N20_25= 30'h3ffe5986,  w8_L2_N20_26= 30'h0007666f,  w8_L2_N20_27= 30'h00013c96,  w8_L2_N20_28= 30'h0004cce1,  w8_L2_N20_29= 30'h3ff969ee;
reg [29:0] w8_L2_N20_30= 30'h00000000,  w8_L2_N20_31= 30'h00038f61,  w8_L2_N20_32= 30'h0009c661,  w8_L2_N20_33= 30'h00000293,  w8_L2_N20_34= 30'h3ffe135f,  w8_L2_N20_35= 30'h0000e172,  w8_L2_N20_36= 30'h3ffffffd,  w8_L2_N20_37= 30'h00000000,  w8_L2_N20_38= 30'h3ffeac2c,  w8_L2_N20_39= 30'h0008c80f,  w8_L2_N20_40= 30'h0001f88c,  w8_L2_N20_41= 30'h3ffdd65b,  w8_L2_N20_42= 30'h00020c95,  w8_L2_N20_43= 30'h00011810,  w8_L2_N20_44= 30'h3ff3c5de,  w8_L2_N20_45= 30'h0002e14c,  w8_L2_N20_46= 30'h0003415a,  w8_L2_N20_47= 30'h3ffd2657,  w8_L2_N20_48= 30'h00000000,  w8_L2_N20_49= 30'h00056400,  w8_L2_N20_50= 30'h00000000,  w8_L2_N20_51= 30'h3fef6d2d,  w8_L2_N20_52= 30'h3ffc9a4c,  w8_L2_N20_53= 30'h0000ebc0,  w8_L2_N20_54= 30'h0001bcd4,  w8_L2_N20_55= 30'h00091d23,  w8_L2_N20_56= 30'h00000003,  w8_L2_N20_57= 30'h00075733,  w8_L2_N20_58= 30'h0007ccef,  w8_L2_N20_59= 30'h0003fa3f;

reg [29:0] w8_out_L_N1_0= 30'h3ffd6f91,  w8_out_L_N1_1= 30'h00000000,  w8_out_L_N1_2= 30'h00006874,  w8_out_L_N1_3= 30'h3fff5ce9,  w8_out_L_N1_4= 30'h000c89d9,  w8_out_L_N1_5= 30'h00000000,  w8_out_L_N1_6= 30'h0009cf4d,  w8_out_L_N1_7= 30'h00000000,  w8_out_L_N1_8= 30'h0003f5af;
reg [29:0] w8_out_L_N1_9= 30'h00000000,  w8_out_L_N1_10= 30'h3ffffb90,  w8_out_L_N1_11= 30'h00000a24,  w8_out_L_N1_12= 30'h00000000,  w8_out_L_N1_13= 30'h00000000,  w8_out_L_N1_14= 30'h0004b34c,  w8_out_L_N1_15= 30'h00000000,  w8_out_L_N1_16= 30'h0002338b,  w8_out_L_N1_17= 30'h3ff75ad2;
reg [29:0] w8_out_L_N1_18= 30'h3ff315d1,  w8_out_L_N1_19= 30'h0008d3b4,  w8_out_L_N2_0= 30'h3ffed834,  w8_out_L_N2_1= 30'h00000000,  w8_out_L_N2_2= 30'h3ff5ea8d,  w8_out_L_N2_3= 30'h0008ad2a,  w8_out_L_N2_4= 30'h000088d6,  w8_out_L_N2_5= 30'h00000000,  w8_out_L_N2_6= 30'h00058d6d;
reg [29:0] w8_out_L_N2_7= 30'h00000000,  w8_out_L_N2_8= 30'h3ff6712d,  w8_out_L_N2_9= 30'h00000000,  w8_out_L_N2_10= 30'h3fff12bb,  w8_out_L_N2_11= 30'h00000000,  w8_out_L_N2_12= 30'h00000000,  w8_out_L_N2_13= 30'h00000000,  w8_out_L_N2_14= 30'h00067e0a,  w8_out_L_N2_15= 30'h00000000;
reg [29:0] w8_out_L_N2_16= 30'h3ff90c1d,  w8_out_L_N2_17= 30'h0008b125,  w8_out_L_N2_18= 30'h3ffa9b57,  w8_out_L_N2_19= 30'h3ffec2db,  w8_out_L_N3_0= 30'h000232fa,  w8_out_L_N3_1= 30'h00000000,  w8_out_L_N3_2= 30'h00035944,  w8_out_L_N3_3= 30'h3fff75be,  w8_out_L_N3_4= 30'h3ff4ca6d;
reg [29:0] w8_out_L_N3_5= 30'h00000000,  w8_out_L_N3_6= 30'h3ff78cec,  w8_out_L_N3_7= 30'h00000000,  w8_out_L_N3_8= 30'h00040c78,  w8_out_L_N3_9= 30'h00000000,  w8_out_L_N3_10= 30'h00008422,  w8_out_L_N3_11= 30'h3fff95eb,  w8_out_L_N3_12= 30'h00000000,  w8_out_L_N3_13= 30'h00000000;
reg [29:0] w8_out_L_N3_14= 30'h3ff37906,  w8_out_L_N3_15= 30'h00000000,  w8_out_L_N3_16= 30'h00050559,  w8_out_L_N3_17= 30'h00006acd,  w8_out_L_N3_18= 30'h000d151a,  w8_out_L_N3_19= 30'h3ffd2c0d; 

reg [58:0] b_L1_N1 = 59'h7ffffee40a561a4,  b_L1_N2 = 59'h7fffff46d1d0eda,  b_L1_N3 = 59'h0000009ce7eb364,  b_L1_N4 = 59'h7fffffef6257a7d,  b_L1_N5 = 59'h7fffff2515a253a,  b_L1_N6 = 59'h7fffff24b702b61,  b_L1_N7 = 59'h7fffffb393d02c0,  b_L1_N8 = 59'h000000f9073a061,  b_L1_N9 = 59'h00000148d8dbced,  b_L1_N10 = 59'h000000c3054dc7b,  b_L1_N11 = 59'h0000013557f432c,  b_L1_N12 = 59'h7fffff73e74afd5,  b_L1_N13 = 59'h0000004a1ba5a2e,  b_L1_N14 = 59'h0000006b296350b,  b_L1_N15 = 59'h00000100b5e6d74,  b_L1_N16 = 59'h7fffff70898e08c,  b_L1_N17 = 59'h7fffffc1c61682d,  b_L1_N18 = 59'h7fffff1dfbf4d88,  b_L1_N19 = 59'h0000003f85c9d90,  b_L1_N20 = 59'h0000009d3600ede,  b_L1_N21 = 59'h000000a5ac7ac7c,  b_L1_N22 = 59'h000001221e2a8d7,  b_L1_N23 = 59'h7fffff4508080c4,  b_L1_N24 = 59'h7ffffefe59dff04,  b_L1_N25 = 59'h000000654481644,  b_L1_N26 = 59'h0000011f4b28477,  b_L1_N27 = 59'h000000ab3bebe97,  b_L1_N28 = 59'h000001af3bfa014,  b_L1_N29 = 59'h0000013d4d19e43,  b_L1_N30 = 59'h0000010d9dd817b;
reg [58:0] b_L1_N31 = 59'h7fffff8f4f3f2d6,  b_L1_N32 = 59'h00000083f6c3c13,  b_L1_N33 = 59'h000000d928f4400,  b_L1_N34 = 59'h7fffff9d115b834,  b_L1_N35 = 59'h0000014506e826a,  b_L1_N36 = 59'h0000012058a6346,  b_L1_N37 = 59'h7fffff0fba780b8,  b_L1_N38 = 59'h7ffffeed6a57e29,  b_L1_N39 = 59'h7fffffc6c2831cd,  b_L1_N40 = 59'h7fffffca499a391,  b_L1_N41 = 59'h000000feac9ad33,  b_L1_N42 = 59'h00000063b83d9ea,  b_L1_N43 = 59'h0000016700022e6,  b_L1_N44 = 59'h0000009a67b9f89,  b_L1_N45 = 59'h0000004ae54400d,  b_L1_N46 = 59'h0000006a2436c10,  b_L1_N47 = 59'h0000010b40ba047,  b_L1_N48 = 59'h0000019f58a0552,  b_L1_N49 = 59'h7fffff3d376d549,  b_L1_N50 = 59'h000000fabefb280,  b_L1_N51 = 59'h7fffff88017dd97,  b_L1_N52 = 59'h000001206c91cea,  b_L1_N53 = 59'h000000902482ec3,  b_L1_N54 = 59'h000000cabb9a1f8,  b_L1_N55 = 59'h000000cdfc4cc22,  b_L1_N56 = 59'h000000a97ee1dd5,  b_L1_N57 = 59'h000000048393c03,  b_L1_N58 = 59'h7fffff7b5e224a3,  b_L1_N59 = 59'h00000095fac62f5,  b_L1_N60 = 59'h000000a3fdac12c;

reg [58:0] b_L2_N1 = 59'h000000df873238e,  b_L2_N2 = 59'h7fffff5aa21f243,  b_L2_N3 = 59'h0000011d84b0537,  b_L2_N4 = 59'h0000009e8abb048,  b_L2_N5 = 59'h000000eb63c11a9,  b_L2_N6 = 59'h7fffff706f78b3c,  b_L2_N7 = 59'h00000069597cc90,  b_L2_N8 = 59'h7fffff198358ba8,  b_L2_N9 = 59'h7fffffa5f1c6566;
reg [58:0] b_L2_N10 = 59'h7fffffc84353f8e,  b_L2_N11 = 59'h00000047d39f79e,  b_L2_N12 = 59'h0000002050cf83f,  b_L2_N13 = 59'h7ffffee7d747faf,  b_L2_N14 = 59'h7fffff852af4f63,  b_L2_N15 = 59'h000000b33a64aad,  b_L2_N16 = 59'h7ffffef7e907ebe,  b_L2_N17 = 59'h0000012a10afd09,  b_L2_N18 = 59'h0000010826aa8eb;
reg [58:0] b_L2_N19 = 59'h7fffffd7dfc7a64,  b_L2_N20 = 59'h7fffff38695050a;

reg [58:0] b_out_L_N1 = 59'h7ffffe94340dcea,  b_out_L_N2 = 59'h7ffffeafba90344,  b_out_L_N3 = 59'h000000b2030acc6;




reg float_a_v;
wire fix_a_v;
reg [31:0]float_a_d;
wire [29:0]fix_a_d;

float_2_fix_6_19 covt_0 ( //32 to 11+19 signed
  .aclk(clk),                                  // input wire aclk
  .s_axis_a_tvalid(float_a_v),            // input wire s_axis_a_tvalid
  .s_axis_a_tdata(float_a_d),              // input wire [31 : 0] s_axis_a_tdata
  .m_axis_result_tvalid(fix_a_v),  // output wire m_axis_result_tvalid
  .m_axis_result_tdata(fix_a_d)    // output wire [23 : 0] m_axis_result_tdata
);


reg [29:0]LBP_161_fix,LBP_156_fix,LBP_137_fix, 
LBP_136_fix,LBP_132_fix,LBP_128_fix,LBP_125_fix,LBP_43_fix,LBP_38_fix,  
LBP_32_fix,LBP_25_fix,LBP_19_fix,LBP_14_fix,LBP_7_fix;

reg [29:0]a_bin198_fix,a_bin199_fix, b_bin208_fix;

reg [29:0]N1_L1=0,N2_L1=0,N3_L1=0,N4_L1=0,N5_L1=0,N6_L1=0,N7_L1=0,N8_L1=0,N9_L1=0,N10_L1=0,
N11_L1=0,N12_L1=0,N13_L1=0,N14_L1=0,N15_L1=0,N16_L1=0,N17_L1=0,N18_L1=0,N19_L1=0,N20_L1=0,N21_L1=0,
N22_L1=0,N23_L1=0,N24_L1=0,N25_L1=0,N26_L1=0,N27_L1=0,N28_L1=0,N29_L1=0,N30_L1=0;
reg [29:0]N31_L1=0,N32_L1=0,N33_L1=0,N34_L1=0,N35_L1=0,N36_L1=0,N37_L1=0,N38_L1=0,N39_L1=0,N40_L1=0,
N41_L1=0,N42_L1=0,N43_L1=0,N44_L1=0,N45_L1=0,N46_L1=0,N47_L1=0,N48_L1=0,N49_L1=0,N50_L1=0,N51_L1=0,
N52_L1=0,N53_L1=0,N54_L1=0,N55_L1=0,N56_L1=0,N57_L1=0,N58_L1=0,N59_L1=0,N60_L1=0;

reg [29:0]N1_L2=0,N2_L2=0,N3_L2=0,N4_L2=0,N5_L2=0,N6_L2=0,N7_L2=0,N8_L2=0,N9_L2=0;
reg [29:0]N10_L2=0,N11_L2=0,N12_L2=0,N13_L2=0,N14_L2=0,N15_L2=0,N16_L2=0,N17_L2=0,N18_L2=0,N19_L2=0,N20_L2=0;

reg [29:0]N1_out_L=0,N2_out_L=0,N3_out_L=0;

localparam [5:0]
st_idle = 0,
st_LBP_161_fix   = 1,
st_LBP_161_fix_s = 2,
st_LBP_156_fix   = 3,
st_LBP_156_fix_s = 4,
st_LBP_137_fix   = 5, 
st_LBP_137_fix_s = 6, 
st_LBP_136_fix   = 7,
st_LBP_136_fix_s = 8,
st_LBP_132_fix   = 9,
st_LBP_132_fix_s = 10,
st_LBP_128_fix   = 11,
st_LBP_128_fix_s = 12,
st_LBP_125_fix   = 13,
st_LBP_125_fix_s = 14,
st_LBP_43_fix    = 15,
st_LBP_43_fix_s  = 16,
st_LBP_38_fix    = 17, 
st_LBP_38_fix_s  = 18,  
st_LBP_32_fix    = 19,
st_LBP_32_fix_s  = 20,
st_LBP_25_fix    = 21,
st_LBP_25_fix_s  = 22,
st_LBP_19_fix    = 23,
st_LBP_19_fix_s  = 24,
st_LBP_14_fix    = 25,
st_LBP_14_fix_s  = 26,
st_LBP_7_fix     = 27,
st_LBP_7_fix_s   = 28,
st_a_bin198_fix  = 29,
st_a_bin198_fix_s= 30,
st_a_bin199_fix  = 31,
st_a_bin199_fix_s= 32,
st_b_bin208_fix  = 33,
st_b_bin208_fix_s= 34,
st_finish        = 35;

reg [5:0]state;
reg fix_done;

always@(posedge clk or posedge reset) 
begin
if(reset)
state <= st_idle;
else
case(state)
    st_idle: begin
    fix_done <= 0;
        if(start_fix_conv) begin
            state <= st_LBP_161_fix;
        end
        else
            state <= st_idle;
    end
    st_LBP_161_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_161;
        state <= st_LBP_161_fix_s;
    end
    st_LBP_161_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_161_fix <= fix_a_d;
            state <= st_LBP_156_fix;
        end   
    end
    st_LBP_156_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_156;
        state <= st_LBP_156_fix_s;
    end
    st_LBP_156_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_156_fix <= fix_a_d;
            state <= st_LBP_137_fix;
        end   
    end
    st_LBP_137_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_137;
        state <= st_LBP_137_fix_s;
    end
    st_LBP_137_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_137_fix <= fix_a_d;
            state <= st_LBP_136_fix;
        end   
    end
    st_LBP_136_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_136;
        state <= st_LBP_136_fix_s;
    end
    st_LBP_136_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_136_fix <= fix_a_d;
            state <= st_LBP_132_fix;
        end   
    end 
    st_LBP_132_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_132;
        state <= st_LBP_132_fix_s;
    end
    st_LBP_132_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_132_fix <= fix_a_d;
            state <= st_LBP_128_fix;
        end   
    end
    st_LBP_128_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_128;
        state <= st_LBP_128_fix_s;
    end
    st_LBP_128_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_128_fix <= fix_a_d;
            state <= st_LBP_125_fix;
        end   
    end
    st_LBP_125_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_125;
        state <= st_LBP_125_fix_s;
    end
    st_LBP_125_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_125_fix <= fix_a_d;
            state <= st_LBP_43_fix;
        end   
    end
    st_LBP_43_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_43;
        state <= st_LBP_43_fix_s;
    end
    st_LBP_43_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_43_fix <= fix_a_d;
            state <= st_LBP_38_fix;
        end   
    end
    st_LBP_38_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_38;
        state <= st_LBP_38_fix_s;
    end
    st_LBP_38_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_38_fix <= fix_a_d;
            state <= st_LBP_32_fix;
        end   
    end
    st_LBP_32_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_32;
        state <= st_LBP_32_fix_s;
    end
    st_LBP_32_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_32_fix <= fix_a_d;
            state <= st_LBP_25_fix;
        end   
    end
    st_LBP_25_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_25;
        state <= st_LBP_25_fix_s;
    end
    st_LBP_25_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_25_fix <= fix_a_d;
            state <= st_LBP_19_fix;
        end   
    end
    st_LBP_19_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_19;
        state <= st_LBP_19_fix_s;
    end
    st_LBP_19_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_19_fix <= fix_a_d;
            state <= st_LBP_14_fix;
        end   
    end
    st_LBP_14_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_14;
        state <= st_LBP_14_fix_s;
    end
    st_LBP_14_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_14_fix <= fix_a_d;
            state <= st_LBP_7_fix;
        end   
    end
    st_LBP_7_fix: begin
        float_a_v <= 1;
        float_a_d <= LBP_7;
        state <= st_LBP_7_fix_s;
    end
    st_LBP_7_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            LBP_7_fix <= fix_a_d;
            state <= st_a_bin198_fix;
        end   
    end
    st_a_bin198_fix: begin
        float_a_v <= 1;
        float_a_d <= a_bin198;
        state <= st_a_bin198_fix_s;
    end
    st_a_bin198_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            a_bin198_fix <= fix_a_d;
            state <= st_a_bin199_fix;
        end   
    end
    st_a_bin199_fix: begin
        float_a_v <= 1;
        float_a_d <= a_bin199;
        state <= st_a_bin199_fix_s;
    end
    st_a_bin199_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            a_bin199_fix <= fix_a_d;
            state <= st_b_bin208_fix;
        end   
    end
    st_b_bin208_fix: begin
        float_a_v <= 1;
        float_a_d <= b_bin208;
        state <= st_b_bin208_fix_s;
    end
    st_b_bin208_fix_s: begin
        float_a_v <= 0;
        if(fix_a_v) begin
            b_bin208_fix <= fix_a_d;
            state <= st_finish;
        end   
    end
    st_finish: begin
        fix_done <= 1;
        state <= st_idle;
    end
    endcase  
end


reg  CE = 0;
reg  [29:0]A,B;
reg  [58:0]C;
wire [58:0]P,PCOUT;
reg  [58:0]NN_aggre;

xbip_multadd_0 your_instance_name (
  .CLK(clk),            // input wire CLK
  .CE(CE),              // input wire CE
  .SCLR(0),          // input wire SCLR
  .A(A),                // input wire [24 : 0] A
  .B(B),                // input wire [24 : 0] B
  .C(C),                // input wire [24 : 0] C
  .SUBTRACT(0),  // input wire SUBTRACT
  .P(P),                // output wire [47 : 0] P
  .PCOUT(PCOUT)        // output wire [47 : 0] PCOUT
);



localparam [5:0]
idle             = 0,
start_L1_NN      = 1,
waiting_L1_NN    = 2,
comp_L1_NN       = 3,    
next_L1_NN       = 4,
done_L1_NN       = 5,
start_L2_NN      = 6,
waiting_L2_NN    = 7,
comp_L2_NN       = 8,
next_L2_NN       = 9,
done_L2_NN       = 10,
start_out_L_NN   = 11,
waiting_out_L_NN = 12,
next_out_L_NN    = 13,
done_out_L_NN    = 14,
compare_outputs  = 15;

reg [5:0]nn_state   = 0;
reg [5:0]count       = 0;
reg [5:0]count_input = 0;
reg [5:0]count_NN    = 0;

always@(posedge clk or posedge reset) 
begin
if(reset) begin
    nn_state    <= idle;
    count       <= 0;
    count_input <= 0;
    NN_aggre    <= 0;
    count_NN    <= 0;
    NN_done     <= 0;
    EB_count    <= 0;
    LB_count    <= 0;
    HD_count    <= 0;
end
else
    case(nn_state)
        idle: begin
                count       <= 0;
                count_input <= 0;
                NN_aggre    <= 0;
                count_NN    <= 0;
                NN_done     <= 0;
            if(fix_done) begin
                nn_state    <= start_L1_NN;
            end else
                nn_state    <= idle;
        end
        start_L1_NN: begin
            case(count_input)
                0: begin
                    A  <= b_bin208_fix; 
                    case(count_NN)
                        0: begin B  <= w8_L1_N1_0;   C  <= b_L1_N1; end
                        1: begin B  <= w8_L1_N2_0;   C  <= b_L1_N2; end
                        2: begin B  <= w8_L1_N3_0;   C  <= b_L1_N3; end
                        3: begin B  <= w8_L1_N4_0;   C  <= b_L1_N4; end
                        4: begin B  <= w8_L1_N5_0;   C  <= b_L1_N5; end
                        5: begin B  <= w8_L1_N6_0;   C  <= b_L1_N6; end
                        6: begin B  <= w8_L1_N7_0;   C  <= b_L1_N7; end
                        7: begin B  <= w8_L1_N8_0;   C  <= b_L1_N8; end
                        8: begin B  <= w8_L1_N9_0;   C  <= b_L1_N9; end
                        9: begin B  <= w8_L1_N10_0;  C  <= b_L1_N10; end
                       10: begin B  <= w8_L1_N11_0;  C  <= b_L1_N11; end
                       11: begin B  <= w8_L1_N12_0;  C  <= b_L1_N12; end
                       12: begin B  <= w8_L1_N13_0;  C  <= b_L1_N13; end
                       13: begin B  <= w8_L1_N14_0;  C  <= b_L1_N14; end
                       14: begin B  <= w8_L1_N15_0;  C  <= b_L1_N15; end
                       15: begin B  <= w8_L1_N16_0;  C  <= b_L1_N16; end
                       16: begin B  <= w8_L1_N17_0;  C  <= b_L1_N17; end
                       17: begin B  <= w8_L1_N18_0;  C  <= b_L1_N18; end
                       18: begin B  <= w8_L1_N19_0;  C  <= b_L1_N19; end
                       19: begin B  <= w8_L1_N20_0;  C  <= b_L1_N20; end
                       20: begin B  <= w8_L1_N21_0;  C  <= b_L1_N21; end
                       21: begin B  <= w8_L1_N22_0;  C  <= b_L1_N22; end
                       22: begin B  <= w8_L1_N23_0;  C  <= b_L1_N23; end
                       23: begin B  <= w8_L1_N24_0;  C  <= b_L1_N24; end
                       24: begin B  <= w8_L1_N25_0;  C  <= b_L1_N25; end
                       25: begin B  <= w8_L1_N26_0;  C  <= b_L1_N26; end
                       26: begin B  <= w8_L1_N27_0;  C  <= b_L1_N27; end
                       27: begin B  <= w8_L1_N28_0;  C  <= b_L1_N28; end
                       28: begin B  <= w8_L1_N29_0;  C  <= b_L1_N29; end
                       29: begin B  <= w8_L1_N30_0;  C  <= b_L1_N30; end
                       30: begin B  <= w8_L1_N31_0;   C  <= b_L1_N31; end
                       31: begin B  <= w8_L1_N32_0;   C  <= b_L1_N32; end
                       32: begin B  <= w8_L1_N33_0;   C  <= b_L1_N33; end
                       33: begin B  <= w8_L1_N34_0;   C  <= b_L1_N34; end
                       34: begin B  <= w8_L1_N35_0;   C  <= b_L1_N35; end
                       35: begin B  <= w8_L1_N36_0;   C  <= b_L1_N36; end
                       36: begin B  <= w8_L1_N37_0;   C  <= b_L1_N37; end
                       37: begin B  <= w8_L1_N38_0;   C  <= b_L1_N38; end
                       38: begin B  <= w8_L1_N39_0;   C  <= b_L1_N39; end
                       39: begin B  <= w8_L1_N40_0;  C  <= b_L1_N40; end
                       40: begin B  <= w8_L1_N41_0;  C  <= b_L1_N41; end
                       41: begin B  <= w8_L1_N42_0;  C  <= b_L1_N42; end
                       42: begin B  <= w8_L1_N43_0;  C  <= b_L1_N43; end
                       43: begin B  <= w8_L1_N44_0;  C  <= b_L1_N44; end
                       44: begin B  <= w8_L1_N45_0;  C  <= b_L1_N45; end
                       45: begin B  <= w8_L1_N46_0;  C  <= b_L1_N46; end
                       46: begin B  <= w8_L1_N47_0;  C  <= b_L1_N47; end
                       47: begin B  <= w8_L1_N48_0;  C  <= b_L1_N48; end
                       48: begin B  <= w8_L1_N49_0;  C  <= b_L1_N49; end
                       49: begin B  <= w8_L1_N50_0;  C  <= b_L1_N50; end
                       50: begin B  <= w8_L1_N51_0;  C  <= b_L1_N51; end
                       51: begin B  <= w8_L1_N52_0;  C  <= b_L1_N52; end
                       52: begin B  <= w8_L1_N53_0;  C  <= b_L1_N53; end
                       53: begin B  <= w8_L1_N54_0;  C  <= b_L1_N54; end
                       54: begin B  <= w8_L1_N55_0;  C  <= b_L1_N55; end
                       55: begin B  <= w8_L1_N56_0;  C  <= b_L1_N56; end
                       56: begin B  <= w8_L1_N57_0;  C  <= b_L1_N57; end
                       57: begin B  <= w8_L1_N58_0;  C  <= b_L1_N58; end
                       58: begin B  <= w8_L1_N59_0;  C  <= b_L1_N59; end
                       59: begin B  <= w8_L1_N60_0;  C  <= b_L1_N60; end
                    endcase
                end
                1: begin
                    A  <= a_bin199_fix; //LBP_161_fix; LBP_156_fix;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_1;
                        1: B  <= w8_L1_N2_1;
                        2: B  <= w8_L1_N3_1;
                        3: B  <= w8_L1_N4_1;
                        4: B  <= w8_L1_N5_1;
                        5: B  <= w8_L1_N6_1;
                        6: B  <= w8_L1_N7_1;
                        7: B  <= w8_L1_N8_1;
                        8: B  <= w8_L1_N9_1;
                        9: B  <= w8_L1_N10_1;
                       10: B  <= w8_L1_N11_1;
                       11: B  <= w8_L1_N12_1;
                       12: B  <= w8_L1_N13_1;
                       13: B  <= w8_L1_N14_1;
                       14: B  <= w8_L1_N15_1;
                       15: B  <= w8_L1_N16_1;
                       16: B  <= w8_L1_N17_1;
                       17: B  <= w8_L1_N18_1;
                       18: B  <= w8_L1_N19_1;
                       19: B  <= w8_L1_N20_1;
                       20: B  <= w8_L1_N21_1;
                       21: B  <= w8_L1_N22_1;
                       22: B  <= w8_L1_N23_1;
                       23: B  <= w8_L1_N24_1;
                       24: B  <= w8_L1_N25_1;
                       25: B  <= w8_L1_N26_1;
                       26: B  <= w8_L1_N27_1;
                       27: B  <= w8_L1_N28_1;
                       28: B  <= w8_L1_N29_1;
                       29: B  <= w8_L1_N30_1;
                       30: B  <= w8_L1_N31_1;
                       31: B  <= w8_L1_N32_1;
                       32: B  <= w8_L1_N33_1;
                       33: B  <= w8_L1_N34_1;
                       34: B  <= w8_L1_N35_1;
                       35: B  <= w8_L1_N36_1;
                       36: B  <= w8_L1_N37_1;
                       37: B  <= w8_L1_N38_1;
                       38: B  <= w8_L1_N39_1;
                       39: B  <= w8_L1_N40_1;
                       40: B  <= w8_L1_N41_1;
                       41: B  <= w8_L1_N42_1;
                       42: B  <= w8_L1_N43_1;
                       43: B  <= w8_L1_N44_1;
                       44: B  <= w8_L1_N45_1;
                       45: B  <= w8_L1_N46_1;
                       46: B  <= w8_L1_N47_1;
                       47: B  <= w8_L1_N48_1;
                       48: B  <= w8_L1_N49_1;
                       49: B  <= w8_L1_N50_1;
                       50: B  <= w8_L1_N51_1;
                       51: B  <= w8_L1_N52_1;
                       52: B  <= w8_L1_N53_1;
                       53: B  <= w8_L1_N54_1;
                       54: B  <= w8_L1_N55_1;
                       55: B  <= w8_L1_N56_1;
                       56: B  <= w8_L1_N57_1;
                       57: B  <= w8_L1_N58_1;
                       58: B  <= w8_L1_N59_1;
                       59: B  <= w8_L1_N60_1;
                    endcase
                end
                2: begin
                    A  <= a_bin198_fix; 
                    B  <= w8_L1_N1_2;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_2;
                        1: B  <= w8_L1_N2_2;
                        2: B  <= w8_L1_N3_2;
                        3: B  <= w8_L1_N4_2;
                        4: B  <= w8_L1_N5_2;
                        5: B  <= w8_L1_N6_2;
                        6: B  <= w8_L1_N7_2;
                        7: B  <= w8_L1_N8_2;
                        8: B  <= w8_L1_N9_2;
                        9: B  <= w8_L1_N10_2;
                       10: B  <= w8_L1_N11_2;
                       11: B  <= w8_L1_N12_2;
                       12: B  <= w8_L1_N13_2;
                       13: B  <= w8_L1_N14_2;
                       14: B  <= w8_L1_N15_2;
                       15: B  <= w8_L1_N16_2;
                       16: B  <= w8_L1_N17_2;
                       17: B  <= w8_L1_N18_2;
                       18: B  <= w8_L1_N19_2;
                       19: B  <= w8_L1_N20_2;
                       20: B  <= w8_L1_N21_2;
                       21: B  <= w8_L1_N22_2;
                       22: B  <= w8_L1_N23_2;
                       23: B  <= w8_L1_N24_2;
                       24: B  <= w8_L1_N25_2;
                       25: B  <= w8_L1_N26_2;
                       26: B  <= w8_L1_N27_2;
                       27: B  <= w8_L1_N28_2;
                       28: B  <= w8_L1_N29_2;
                       29: B  <= w8_L1_N30_2;
                       30: B  <= w8_L1_N31_2;
                       31: B  <= w8_L1_N32_2;
                       32: B  <= w8_L1_N33_2;
                       33: B  <= w8_L1_N34_2;
                       34: B  <= w8_L1_N35_2;
                       35: B  <= w8_L1_N36_2;
                       36: B  <= w8_L1_N37_2;
                       37: B  <= w8_L1_N38_2;
                       38: B  <= w8_L1_N39_2;
                       39: B  <= w8_L1_N40_2;
                       40: B  <= w8_L1_N41_2;
                       41: B  <= w8_L1_N42_2;
                       42: B  <= w8_L1_N43_2;
                       43: B  <= w8_L1_N44_2;
                       44: B  <= w8_L1_N45_2;
                       45: B  <= w8_L1_N46_2;
                       46: B  <= w8_L1_N47_2;
                       47: B  <= w8_L1_N48_2;
                       48: B  <= w8_L1_N49_2;
                       49: B  <= w8_L1_N50_2;
                       50: B  <= w8_L1_N51_2;
                       51: B  <= w8_L1_N52_2;
                       52: B  <= w8_L1_N53_2;
                       53: B  <= w8_L1_N54_2;
                       54: B  <= w8_L1_N55_2;
                       55: B  <= w8_L1_N56_2;
                       56: B  <= w8_L1_N57_2;
                       57: B  <= w8_L1_N58_2;
                       58: B  <= w8_L1_N59_2;
                       59: B  <= w8_L1_N60_2;
                    endcase
                end
                3: begin
                    A  <= LBP_161_fix; //LBP_161
                    B  <= w8_L1_N1_3;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_3;
                        1: B  <= w8_L1_N2_3;
                        2: B  <= w8_L1_N3_3;
                        3: B  <= w8_L1_N4_3;
                        4: B  <= w8_L1_N5_3;
                        5: B  <= w8_L1_N6_3;
                        6: B  <= w8_L1_N7_3;
                        7: B  <= w8_L1_N8_3;
                        8: B  <= w8_L1_N9_3;
                        9: B  <= w8_L1_N10_3;
                       10: B  <= w8_L1_N11_3;
                       11: B  <= w8_L1_N12_3;
                       12: B  <= w8_L1_N13_3;
                       13: B  <= w8_L1_N14_3;
                       14: B  <= w8_L1_N15_3;
                       15: B  <= w8_L1_N16_3;
                       16: B  <= w8_L1_N17_3;
                       17: B  <= w8_L1_N18_3;
                       18: B  <= w8_L1_N19_3;
                       19: B  <= w8_L1_N20_3;
                       20: B  <= w8_L1_N21_3;
                       21: B  <= w8_L1_N22_3;
                       22: B  <= w8_L1_N23_3;
                       23: B  <= w8_L1_N24_3;
                       24: B  <= w8_L1_N25_3;
                       25: B  <= w8_L1_N26_3;
                       26: B  <= w8_L1_N27_3;
                       27: B  <= w8_L1_N28_3;
                       28: B  <= w8_L1_N29_3;
                       29: B  <= w8_L1_N30_3;
                       30: B  <= w8_L1_N31_3;
                       31: B  <= w8_L1_N32_3;
                       32: B  <= w8_L1_N33_3;
                       33: B  <= w8_L1_N34_3;
                       34: B  <= w8_L1_N35_3;
                       35: B  <= w8_L1_N36_3;
                       36: B  <= w8_L1_N37_3;
                       37: B  <= w8_L1_N38_3;
                       38: B  <= w8_L1_N39_3;
                       39: B  <= w8_L1_N40_3;
                       40: B  <= w8_L1_N41_3;
                       41: B  <= w8_L1_N42_3;
                       42: B  <= w8_L1_N43_3;
                       43: B  <= w8_L1_N44_3;
                       44: B  <= w8_L1_N45_3;
                       45: B  <= w8_L1_N46_3;
                       46: B  <= w8_L1_N47_3;
                       47: B  <= w8_L1_N48_3;
                       48: B  <= w8_L1_N49_3;
                       49: B  <= w8_L1_N50_3;
                       50: B  <= w8_L1_N51_3;
                       51: B  <= w8_L1_N52_3;
                       52: B  <= w8_L1_N53_3;
                       53: B  <= w8_L1_N54_3;
                       54: B  <= w8_L1_N55_3;
                       55: B  <= w8_L1_N56_3;
                       56: B  <= w8_L1_N57_3;
                       57: B  <= w8_L1_N58_3;
                       58: B  <= w8_L1_N59_3;
                       59: B  <= w8_L1_N60_3;
                    endcase
                end
                4: begin
                    A  <= LBP_156_fix; 
                    B  <= w8_L1_N1_4;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_4;
                        1: B  <= w8_L1_N2_4;
                        2: B  <= w8_L1_N3_4;
                        3: B  <= w8_L1_N4_4;
                        4: B  <= w8_L1_N5_4;
                        5: B  <= w8_L1_N6_4;
                        6: B  <= w8_L1_N7_4;
                        7: B  <= w8_L1_N8_4;
                        8: B  <= w8_L1_N9_4;
                        9: B  <= w8_L1_N10_4;
                       10: B  <= w8_L1_N11_4;
                       11: B  <= w8_L1_N12_4;
                       12: B  <= w8_L1_N13_4;
                       13: B  <= w8_L1_N14_4;
                       14: B  <= w8_L1_N15_4;
                       15: B  <= w8_L1_N16_4;
                       16: B  <= w8_L1_N17_4;
                       17: B  <= w8_L1_N18_4;
                       18: B  <= w8_L1_N19_4;
                       19: B  <= w8_L1_N20_4;
                       20: B  <= w8_L1_N21_4;
                       21: B  <= w8_L1_N22_4;
                       22: B  <= w8_L1_N23_4;
                       23: B  <= w8_L1_N24_4;
                       24: B  <= w8_L1_N25_4;
                       25: B  <= w8_L1_N26_4;
                       26: B  <= w8_L1_N27_4;
                       27: B  <= w8_L1_N28_4;
                       28: B  <= w8_L1_N29_4;
                       29: B  <= w8_L1_N30_4;
                       30: B  <= w8_L1_N31_4;
                       31: B  <= w8_L1_N32_4;
                       32: B  <= w8_L1_N33_4;
                       33: B  <= w8_L1_N34_4;
                       34: B  <= w8_L1_N35_4;
                       35: B  <= w8_L1_N36_4;
                       36: B  <= w8_L1_N37_4;
                       37: B  <= w8_L1_N38_4;
                       38: B  <= w8_L1_N39_4;
                       39: B  <= w8_L1_N40_4;
                       40: B  <= w8_L1_N41_4;
                       41: B  <= w8_L1_N42_4;
                       42: B  <= w8_L1_N43_4;
                       43: B  <= w8_L1_N44_4;
                       44: B  <= w8_L1_N45_4;
                       45: B  <= w8_L1_N46_4;
                       46: B  <= w8_L1_N47_4;
                       47: B  <= w8_L1_N48_4;
                       48: B  <= w8_L1_N49_4;
                       49: B  <= w8_L1_N50_4;
                       50: B  <= w8_L1_N51_4;
                       51: B  <= w8_L1_N52_4;
                       52: B  <= w8_L1_N53_4;
                       53: B  <= w8_L1_N54_4;
                       54: B  <= w8_L1_N55_4;
                       55: B  <= w8_L1_N56_4;
                       56: B  <= w8_L1_N57_4;
                       57: B  <= w8_L1_N58_4;
                       58: B  <= w8_L1_N59_4;
                       59: B  <= w8_L1_N60_4;
                    endcase
                end
                5: begin
                    A  <= LBP_137_fix;
                    B  <= w8_L1_N1_5;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_5;
                        1: B  <= w8_L1_N2_5;
                        2: B  <= w8_L1_N3_5;
                        3: B  <= w8_L1_N4_5;
                        4: B  <= w8_L1_N5_5;
                        5: B  <= w8_L1_N6_5;
                        6: B  <= w8_L1_N7_5;
                        7: B  <= w8_L1_N8_5;
                        8: B  <= w8_L1_N9_5;
                        9: B  <= w8_L1_N10_5;
                       10: B  <= w8_L1_N11_5;
                       11: B  <= w8_L1_N12_5;
                       12: B  <= w8_L1_N13_5;
                       13: B  <= w8_L1_N14_5;
                       14: B  <= w8_L1_N15_5;
                       15: B  <= w8_L1_N16_5;
                       16: B  <= w8_L1_N17_5;
                       17: B  <= w8_L1_N18_5;
                       18: B  <= w8_L1_N19_5;
                       19: B  <= w8_L1_N20_5;
                       20: B  <= w8_L1_N21_5;
                       21: B  <= w8_L1_N22_5;
                       22: B  <= w8_L1_N23_5;
                       23: B  <= w8_L1_N24_5;
                       24: B  <= w8_L1_N25_5;
                       25: B  <= w8_L1_N26_5;
                       26: B  <= w8_L1_N27_5;
                       27: B  <= w8_L1_N28_5;
                       28: B  <= w8_L1_N29_5;
                       29: B  <= w8_L1_N30_5;
                       30: B  <= w8_L1_N31_5;
                       31: B  <= w8_L1_N32_5;
                       32: B  <= w8_L1_N33_5;
                       33: B  <= w8_L1_N34_5;
                       34: B  <= w8_L1_N35_5;
                       35: B  <= w8_L1_N36_5;
                       36: B  <= w8_L1_N37_5;
                       37: B  <= w8_L1_N38_5;
                       38: B  <= w8_L1_N39_5;
                       39: B  <= w8_L1_N40_5;
                       40: B  <= w8_L1_N41_5;
                       41: B  <= w8_L1_N42_5;
                       42: B  <= w8_L1_N43_5;
                       43: B  <= w8_L1_N44_5;
                       44: B  <= w8_L1_N45_5;
                       45: B  <= w8_L1_N46_5;
                       46: B  <= w8_L1_N47_5;
                       47: B  <= w8_L1_N48_5;
                       48: B  <= w8_L1_N49_5;
                       49: B  <= w8_L1_N50_5;
                       50: B  <= w8_L1_N51_5;
                       51: B  <= w8_L1_N52_5;
                       52: B  <= w8_L1_N53_5;
                       53: B  <= w8_L1_N54_5;
                       54: B  <= w8_L1_N55_5;
                       55: B  <= w8_L1_N56_5;
                       56: B  <= w8_L1_N57_5;
                       57: B  <= w8_L1_N58_5;
                       58: B  <= w8_L1_N59_5;
                       59: B  <= w8_L1_N60_5;
                    endcase
                end
                6: begin
                    A  <= LBP_136_fix;
                    B  <= w8_L1_N1_6;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_6;
                        1: B  <= w8_L1_N2_6;
                        2: B  <= w8_L1_N3_6;
                        3: B  <= w8_L1_N4_6;
                        4: B  <= w8_L1_N5_6;
                        5: B  <= w8_L1_N6_6;
                        6: B  <= w8_L1_N7_6;
                        7: B  <= w8_L1_N8_6;
                        8: B  <= w8_L1_N9_6;
                        9: B  <= w8_L1_N10_6;
                       10: B  <= w8_L1_N11_6;
                       11: B  <= w8_L1_N12_6;
                       12: B  <= w8_L1_N13_6;
                       13: B  <= w8_L1_N14_6;
                       14: B  <= w8_L1_N15_6;
                       15: B  <= w8_L1_N16_6;
                       16: B  <= w8_L1_N17_6;
                       17: B  <= w8_L1_N18_6;
                       18: B  <= w8_L1_N19_6;
                       19: B  <= w8_L1_N20_6;
                       20: B  <= w8_L1_N21_6;
                       21: B  <= w8_L1_N22_6;
                       22: B  <= w8_L1_N23_6;
                       23: B  <= w8_L1_N24_6;
                       24: B  <= w8_L1_N25_6;
                       25: B  <= w8_L1_N26_6;
                       26: B  <= w8_L1_N27_6;
                       27: B  <= w8_L1_N28_6;
                       28: B  <= w8_L1_N29_6;
                       29: B  <= w8_L1_N30_6;
                       30: B  <= w8_L1_N31_6;
                       31: B  <= w8_L1_N32_6;
                       32: B  <= w8_L1_N33_6;
                       33: B  <= w8_L1_N34_6;
                       34: B  <= w8_L1_N35_6;
                       35: B  <= w8_L1_N36_6;
                       36: B  <= w8_L1_N37_6;
                       37: B  <= w8_L1_N38_6;
                       38: B  <= w8_L1_N39_6;
                       39: B  <= w8_L1_N40_6;
                       40: B  <= w8_L1_N41_6;
                       41: B  <= w8_L1_N42_6;
                       42: B  <= w8_L1_N43_6;
                       43: B  <= w8_L1_N44_6;
                       44: B  <= w8_L1_N45_6;
                       45: B  <= w8_L1_N46_6;
                       46: B  <= w8_L1_N47_6;
                       47: B  <= w8_L1_N48_6;
                       48: B  <= w8_L1_N49_6;
                       49: B  <= w8_L1_N50_6;
                       50: B  <= w8_L1_N51_6;
                       51: B  <= w8_L1_N52_6;
                       52: B  <= w8_L1_N53_6;
                       53: B  <= w8_L1_N54_6;
                       54: B  <= w8_L1_N55_6;
                       55: B  <= w8_L1_N56_6;
                       56: B  <= w8_L1_N57_6;
                       57: B  <= w8_L1_N58_6;
                       58: B  <= w8_L1_N59_6;
                       59: B  <= w8_L1_N60_6;
                    endcase
                end
                7: begin
                    A  <= LBP_132_fix;     
                    B  <= w8_L1_N1_7;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_7;
                        1: B  <= w8_L1_N2_7;
                        2: B  <= w8_L1_N3_7;
                        3: B  <= w8_L1_N4_7;
                        4: B  <= w8_L1_N5_7;
                        5: B  <= w8_L1_N6_7;
                        6: B  <= w8_L1_N7_7;
                        7: B  <= w8_L1_N8_7;
                        8: B  <= w8_L1_N9_7;
                        9: B  <= w8_L1_N10_7;
                       10: B  <= w8_L1_N11_7;
                       11: B  <= w8_L1_N12_7;
                       12: B  <= w8_L1_N13_7;
                       13: B  <= w8_L1_N14_7;
                       14: B  <= w8_L1_N15_7;
                       15: B  <= w8_L1_N16_7;
                       16: B  <= w8_L1_N17_7;
                       17: B  <= w8_L1_N18_7;
                       18: B  <= w8_L1_N19_7;
                       19: B  <= w8_L1_N20_7;
                       20: B  <= w8_L1_N21_7;
                       21: B  <= w8_L1_N22_7;
                       22: B  <= w8_L1_N23_7;
                       23: B  <= w8_L1_N24_7;
                       24: B  <= w8_L1_N25_7;
                       25: B  <= w8_L1_N26_7;
                       26: B  <= w8_L1_N27_7;
                       27: B  <= w8_L1_N28_7;
                       28: B  <= w8_L1_N29_7;
                       29: B  <= w8_L1_N30_7;
                       30: B  <= w8_L1_N31_7;
                       31: B  <= w8_L1_N32_7;
                       32: B  <= w8_L1_N33_7;
                       33: B  <= w8_L1_N34_7;
                       34: B  <= w8_L1_N35_7;
                       35: B  <= w8_L1_N36_7;
                       36: B  <= w8_L1_N37_7;
                       37: B  <= w8_L1_N38_7;
                       38: B  <= w8_L1_N39_7;
                       39: B  <= w8_L1_N40_7;
                       40: B  <= w8_L1_N41_7;
                       41: B  <= w8_L1_N42_7;
                       42: B  <= w8_L1_N43_7;
                       43: B  <= w8_L1_N44_7;
                       44: B  <= w8_L1_N45_7;
                       45: B  <= w8_L1_N46_7;
                       46: B  <= w8_L1_N47_7;
                       47: B  <= w8_L1_N48_7;
                       48: B  <= w8_L1_N49_7;
                       49: B  <= w8_L1_N50_7;
                       50: B  <= w8_L1_N51_7;
                       51: B  <= w8_L1_N52_7;
                       52: B  <= w8_L1_N53_7;
                       53: B  <= w8_L1_N54_7;
                       54: B  <= w8_L1_N55_7;
                       55: B  <= w8_L1_N56_7;
                       56: B  <= w8_L1_N57_7;
                       57: B  <= w8_L1_N58_7;
                       58: B  <= w8_L1_N59_7;
                       59: B  <= w8_L1_N60_7;
                    endcase
                end
                8: begin
                    A  <= LBP_128_fix;  
                    B  <= w8_L1_N1_8;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_8;
                        1: B  <= w8_L1_N2_8;
                        2: B  <= w8_L1_N3_8;
                        3: B  <= w8_L1_N4_8;
                        4: B  <= w8_L1_N5_8;
                        5: B  <= w8_L1_N6_8;
                        6: B  <= w8_L1_N7_8;
                        7: B  <= w8_L1_N8_8;
                        8: B  <= w8_L1_N9_8;
                        9: B  <= w8_L1_N10_8;
                       10: B  <= w8_L1_N11_8;
                       11: B  <= w8_L1_N12_8;
                       12: B  <= w8_L1_N13_8;
                       13: B  <= w8_L1_N14_8;
                       14: B  <= w8_L1_N15_8;
                       15: B  <= w8_L1_N16_8;
                       16: B  <= w8_L1_N17_8;
                       17: B  <= w8_L1_N18_8;
                       18: B  <= w8_L1_N19_8;
                       19: B  <= w8_L1_N20_8;
                       20: B  <= w8_L1_N21_8;
                       21: B  <= w8_L1_N22_8;
                       22: B  <= w8_L1_N23_8;
                       23: B  <= w8_L1_N24_8;
                       24: B  <= w8_L1_N25_8;
                       25: B  <= w8_L1_N26_8;
                       26: B  <= w8_L1_N27_8;
                       27: B  <= w8_L1_N28_8;
                       28: B  <= w8_L1_N29_8;
                       29: B  <= w8_L1_N30_8;
                       30: B  <= w8_L1_N31_8;
                       31: B  <= w8_L1_N32_8;
                       32: B  <= w8_L1_N33_8;
                       33: B  <= w8_L1_N34_8;
                       34: B  <= w8_L1_N35_8;
                       35: B  <= w8_L1_N36_8;
                       36: B  <= w8_L1_N37_8;
                       37: B  <= w8_L1_N38_8;
                       38: B  <= w8_L1_N39_8;
                       39: B  <= w8_L1_N40_8;
                       40: B  <= w8_L1_N41_8;
                       41: B  <= w8_L1_N42_8;
                       42: B  <= w8_L1_N43_8;
                       43: B  <= w8_L1_N44_8;
                       44: B  <= w8_L1_N45_8;
                       45: B  <= w8_L1_N46_8;
                       46: B  <= w8_L1_N47_8;
                       47: B  <= w8_L1_N48_8;
                       48: B  <= w8_L1_N49_8;
                       49: B  <= w8_L1_N50_8;
                       50: B  <= w8_L1_N51_8;
                       51: B  <= w8_L1_N52_8;
                       52: B  <= w8_L1_N53_8;
                       53: B  <= w8_L1_N54_8;
                       54: B  <= w8_L1_N55_8;
                       55: B  <= w8_L1_N56_8;
                       56: B  <= w8_L1_N57_8;
                       57: B  <= w8_L1_N58_8;
                       58: B  <= w8_L1_N59_8;
                       59: B  <= w8_L1_N60_8;
                    endcase
                end
                9: begin
                    A  <= LBP_125_fix;
                    B  <= w8_L1_N1_9;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_9;
                        1: B  <= w8_L1_N2_9;
                        2: B  <= w8_L1_N3_9;
                        3: B  <= w8_L1_N4_9;
                        4: B  <= w8_L1_N5_9;
                        5: B  <= w8_L1_N6_9;
                        6: B  <= w8_L1_N7_9;
                        7: B  <= w8_L1_N8_9;
                        8: B  <= w8_L1_N9_9;
                        9: B  <= w8_L1_N10_9;
                       10: B  <= w8_L1_N11_9;
                       11: B  <= w8_L1_N12_9;
                       12: B  <= w8_L1_N13_9;
                       13: B  <= w8_L1_N14_9;
                       14: B  <= w8_L1_N15_9;
                       15: B  <= w8_L1_N16_9;
                       16: B  <= w8_L1_N17_9;
                       17: B  <= w8_L1_N18_9;
                       18: B  <= w8_L1_N19_9;
                       19: B  <= w8_L1_N20_9;
                       20: B  <= w8_L1_N21_9;
                       21: B  <= w8_L1_N22_9;
                       22: B  <= w8_L1_N23_9;
                       23: B  <= w8_L1_N24_9;
                       24: B  <= w8_L1_N25_9;
                       25: B  <= w8_L1_N26_9;
                       26: B  <= w8_L1_N27_9;
                       27: B  <= w8_L1_N28_9;
                       28: B  <= w8_L1_N29_9;
                       29: B  <= w8_L1_N30_9;
                       30: B  <= w8_L1_N31_9;
                       31: B  <= w8_L1_N32_9;
                       32: B  <= w8_L1_N33_9;
                       33: B  <= w8_L1_N34_9;
                       34: B  <= w8_L1_N35_9;
                       35: B  <= w8_L1_N36_9;
                       36: B  <= w8_L1_N37_9;
                       37: B  <= w8_L1_N38_9;
                       38: B  <= w8_L1_N39_9;
                       39: B  <= w8_L1_N40_9;
                       40: B  <= w8_L1_N41_9;
                       41: B  <= w8_L1_N42_9;
                       42: B  <= w8_L1_N43_9;
                       43: B  <= w8_L1_N44_9;
                       44: B  <= w8_L1_N45_9;
                       45: B  <= w8_L1_N46_9;
                       46: B  <= w8_L1_N47_9;
                       47: B  <= w8_L1_N48_9;
                       48: B  <= w8_L1_N49_9;
                       49: B  <= w8_L1_N50_9;
                       50: B  <= w8_L1_N51_9;
                       51: B  <= w8_L1_N52_9;
                       52: B  <= w8_L1_N53_9;
                       53: B  <= w8_L1_N54_9;
                       54: B  <= w8_L1_N55_9;
                       55: B  <= w8_L1_N56_9;
                       56: B  <= w8_L1_N57_9;
                       57: B  <= w8_L1_N58_9;
                       58: B  <= w8_L1_N59_9;
                       59: B  <= w8_L1_N60_9;
                    endcase
                end
                10: begin
                    A  <= LBP_43_fix;    
                    B  <= w8_L1_N1_10;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_10;
                        1: B  <= w8_L1_N2_10;
                        2: B  <= w8_L1_N3_10;
                        3: B  <= w8_L1_N4_10;
                        4: B  <= w8_L1_N5_10;
                        5: B  <= w8_L1_N6_10;
                        6: B  <= w8_L1_N7_10;
                        7: B  <= w8_L1_N8_10;
                        8: B  <= w8_L1_N9_10;
                        9: B  <= w8_L1_N10_10;
                       10: B  <= w8_L1_N11_10;
                       11: B  <= w8_L1_N12_10;
                       12: B  <= w8_L1_N13_10;
                       13: B  <= w8_L1_N14_10;
                       14: B  <= w8_L1_N15_10;
                       15: B  <= w8_L1_N16_10;
                       16: B  <= w8_L1_N17_10;
                       17: B  <= w8_L1_N18_10;
                       18: B  <= w8_L1_N19_10;
                       19: B  <= w8_L1_N20_10;
                       20: B  <= w8_L1_N21_10;
                       21: B  <= w8_L1_N22_10;
                       22: B  <= w8_L1_N23_10;
                       23: B  <= w8_L1_N24_10;
                       24: B  <= w8_L1_N25_10;
                       25: B  <= w8_L1_N26_10;
                       26: B  <= w8_L1_N27_10;
                       27: B  <= w8_L1_N28_10;
                       28: B  <= w8_L1_N29_10;
                       29: B  <= w8_L1_N30_10;
                       30: B  <= w8_L1_N31_10;
                       31: B  <= w8_L1_N32_10;
                       32: B  <= w8_L1_N33_10;
                       33: B  <= w8_L1_N34_10;
                       34: B  <= w8_L1_N35_10;
                       35: B  <= w8_L1_N36_10;
                       36: B  <= w8_L1_N37_10;
                       37: B  <= w8_L1_N38_10;
                       38: B  <= w8_L1_N39_10;
                       39: B  <= w8_L1_N40_10;
                       40: B  <= w8_L1_N41_10;
                       41: B  <= w8_L1_N42_10;
                       42: B  <= w8_L1_N43_10;
                       43: B  <= w8_L1_N44_10;
                       44: B  <= w8_L1_N45_10;
                       45: B  <= w8_L1_N46_10;
                       46: B  <= w8_L1_N47_10;
                       47: B  <= w8_L1_N48_10;
                       48: B  <= w8_L1_N49_10;
                       49: B  <= w8_L1_N50_10;
                       50: B  <= w8_L1_N51_10;
                       51: B  <= w8_L1_N52_10;
                       52: B  <= w8_L1_N53_10;
                       53: B  <= w8_L1_N54_10;
                       54: B  <= w8_L1_N55_10;
                       55: B  <= w8_L1_N56_10;
                       56: B  <= w8_L1_N57_10;
                       57: B  <= w8_L1_N58_10;
                       58: B  <= w8_L1_N59_10;
                       59: B  <= w8_L1_N60_10;
                    endcase
                end
                11: begin
                    A  <= LBP_38_fix;   
                    B  <= w8_L1_N1_11;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_11;
                        1: B  <= w8_L1_N2_11;
                        2: B  <= w8_L1_N3_11;
                        3: B  <= w8_L1_N4_11;
                        4: B  <= w8_L1_N5_11;
                        5: B  <= w8_L1_N6_11;
                        6: B  <= w8_L1_N7_11;
                        7: B  <= w8_L1_N8_11;
                        8: B  <= w8_L1_N9_11;
                        9: B  <= w8_L1_N10_11;
                       10: B  <= w8_L1_N11_11;
                       11: B  <= w8_L1_N12_11;
                       12: B  <= w8_L1_N13_11;
                       13: B  <= w8_L1_N14_11;
                       14: B  <= w8_L1_N15_11;
                       15: B  <= w8_L1_N16_11;
                       16: B  <= w8_L1_N17_11;
                       17: B  <= w8_L1_N18_11;
                       18: B  <= w8_L1_N19_11;
                       19: B  <= w8_L1_N20_11;
                       20: B  <= w8_L1_N21_11;
                       21: B  <= w8_L1_N22_11;
                       22: B  <= w8_L1_N23_11;
                       23: B  <= w8_L1_N24_11;
                       24: B  <= w8_L1_N25_11;
                       25: B  <= w8_L1_N26_11;
                       26: B  <= w8_L1_N27_11;
                       27: B  <= w8_L1_N28_11;
                       28: B  <= w8_L1_N29_11;
                       29: B  <= w8_L1_N30_11;
                       30: B  <= w8_L1_N31_11;
                       31: B  <= w8_L1_N32_11;
                       32: B  <= w8_L1_N33_11;
                       33: B  <= w8_L1_N34_11;
                       34: B  <= w8_L1_N35_11;
                       35: B  <= w8_L1_N36_11;
                       36: B  <= w8_L1_N37_11;
                       37: B  <= w8_L1_N38_11;
                       38: B  <= w8_L1_N39_11;
                       39: B  <= w8_L1_N40_11;
                       40: B  <= w8_L1_N41_11;
                       41: B  <= w8_L1_N42_11;
                       42: B  <= w8_L1_N43_11;
                       43: B  <= w8_L1_N44_11;
                       44: B  <= w8_L1_N45_11;
                       45: B  <= w8_L1_N46_11;
                       46: B  <= w8_L1_N47_11;
                       47: B  <= w8_L1_N48_11;
                       48: B  <= w8_L1_N49_11;
                       49: B  <= w8_L1_N50_11;
                       50: B  <= w8_L1_N51_11;
                       51: B  <= w8_L1_N52_11;
                       52: B  <= w8_L1_N53_11;
                       53: B  <= w8_L1_N54_11;
                       54: B  <= w8_L1_N55_11;
                       55: B  <= w8_L1_N56_11;
                       56: B  <= w8_L1_N57_11;
                       57: B  <= w8_L1_N58_11;
                       58: B  <= w8_L1_N59_11;
                       59: B  <= w8_L1_N60_11;
                    endcase
                end
                12: begin
                    A  <= LBP_32_fix;    
                    B  <= w8_L1_N1_12;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_12;
                        1: B  <= w8_L1_N2_12;
                        2: B  <= w8_L1_N3_12;
                        3: B  <= w8_L1_N4_12;
                        4: B  <= w8_L1_N5_12;
                        5: B  <= w8_L1_N6_12;
                        6: B  <= w8_L1_N7_12;
                        7: B  <= w8_L1_N8_12;
                        8: B  <= w8_L1_N9_12;
                        9: B  <= w8_L1_N10_12;
                       10: B  <= w8_L1_N11_12;
                       11: B  <= w8_L1_N12_12;
                       12: B  <= w8_L1_N13_12;
                       13: B  <= w8_L1_N14_12;
                       14: B  <= w8_L1_N15_12;
                       15: B  <= w8_L1_N16_12;
                       16: B  <= w8_L1_N17_12;
                       17: B  <= w8_L1_N18_12;
                       18: B  <= w8_L1_N19_12;
                       19: B  <= w8_L1_N20_12;
                       20: B  <= w8_L1_N21_12;
                       21: B  <= w8_L1_N22_12;
                       22: B  <= w8_L1_N23_12;
                       23: B  <= w8_L1_N24_12;
                       24: B  <= w8_L1_N25_12;
                       25: B  <= w8_L1_N26_12;
                       26: B  <= w8_L1_N27_12;
                       27: B  <= w8_L1_N28_12;
                       28: B  <= w8_L1_N29_12;
                       29: B  <= w8_L1_N30_12;
                       30: B  <= w8_L1_N31_12;
                       31: B  <= w8_L1_N32_12;
                       32: B  <= w8_L1_N33_12;
                       33: B  <= w8_L1_N34_12;
                       34: B  <= w8_L1_N35_12;
                       35: B  <= w8_L1_N36_12;
                       36: B  <= w8_L1_N37_12;
                       37: B  <= w8_L1_N38_12;
                       38: B  <= w8_L1_N39_12;
                       39: B  <= w8_L1_N40_12;
                       40: B  <= w8_L1_N41_12;
                       41: B  <= w8_L1_N42_12;
                       42: B  <= w8_L1_N43_12;
                       43: B  <= w8_L1_N44_12;
                       44: B  <= w8_L1_N45_12;
                       45: B  <= w8_L1_N46_12;
                       46: B  <= w8_L1_N47_12;
                       47: B  <= w8_L1_N48_12;
                       48: B  <= w8_L1_N49_12;
                       49: B  <= w8_L1_N50_12;
                       50: B  <= w8_L1_N51_12;
                       51: B  <= w8_L1_N52_12;
                       52: B  <= w8_L1_N53_12;
                       53: B  <= w8_L1_N54_12;
                       54: B  <= w8_L1_N55_12;
                       55: B  <= w8_L1_N56_12;
                       56: B  <= w8_L1_N57_12;
                       57: B  <= w8_L1_N58_12;
                       58: B  <= w8_L1_N59_12;
                       59: B  <= w8_L1_N60_12;
                    endcase
                end
                13: begin
                    A  <= LBP_25_fix;   
                    B  <= w8_L1_N1_13;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_13;
                        1: B  <= w8_L1_N2_13;
                        2: B  <= w8_L1_N3_13;
                        3: B  <= w8_L1_N4_13;
                        4: B  <= w8_L1_N5_13;
                        5: B  <= w8_L1_N6_13;
                        6: B  <= w8_L1_N7_13;
                        7: B  <= w8_L1_N8_13;
                        8: B  <= w8_L1_N9_13;
                        9: B  <= w8_L1_N10_13;
                       10: B  <= w8_L1_N11_13;
                       11: B  <= w8_L1_N12_13;
                       12: B  <= w8_L1_N13_13;
                       13: B  <= w8_L1_N14_13;
                       14: B  <= w8_L1_N15_13;
                       15: B  <= w8_L1_N16_13;
                       16: B  <= w8_L1_N17_13;
                       17: B  <= w8_L1_N18_13;
                       18: B  <= w8_L1_N19_13;
                       19: B  <= w8_L1_N20_13;
                       20: B  <= w8_L1_N21_13;
                       21: B  <= w8_L1_N22_13;
                       22: B  <= w8_L1_N23_13;
                       23: B  <= w8_L1_N24_13;
                       24: B  <= w8_L1_N25_13;
                       25: B  <= w8_L1_N26_13;
                       26: B  <= w8_L1_N27_13;
                       27: B  <= w8_L1_N28_13;
                       28: B  <= w8_L1_N29_13;
                       29: B  <= w8_L1_N30_13;
                       30: B  <= w8_L1_N31_13;
                       31: B  <= w8_L1_N32_13;
                       32: B  <= w8_L1_N33_13;
                       33: B  <= w8_L1_N34_13;
                       34: B  <= w8_L1_N35_13;
                       35: B  <= w8_L1_N36_13;
                       36: B  <= w8_L1_N37_13;
                       37: B  <= w8_L1_N38_13;
                       38: B  <= w8_L1_N39_13;
                       39: B  <= w8_L1_N40_13;
                       40: B  <= w8_L1_N41_13;
                       41: B  <= w8_L1_N42_13;
                       42: B  <= w8_L1_N43_13;
                       43: B  <= w8_L1_N44_13;
                       44: B  <= w8_L1_N45_13;
                       45: B  <= w8_L1_N46_13;
                       46: B  <= w8_L1_N47_13;
                       47: B  <= w8_L1_N48_13;
                       48: B  <= w8_L1_N49_13;
                       49: B  <= w8_L1_N50_13;
                       50: B  <= w8_L1_N51_13;
                       51: B  <= w8_L1_N52_13;
                       52: B  <= w8_L1_N53_13;
                       53: B  <= w8_L1_N54_13;
                       54: B  <= w8_L1_N55_13;
                       55: B  <= w8_L1_N56_13;
                       56: B  <= w8_L1_N57_13;
                       57: B  <= w8_L1_N58_13;
                       58: B  <= w8_L1_N59_13;
                       59: B  <= w8_L1_N60_13;
                    endcase
                end
                14: begin
                    A  <= LBP_19_fix;  
                    B  <= w8_L1_N1_14;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_14;
                        1: B  <= w8_L1_N2_14;
                        2: B  <= w8_L1_N3_14;
                        3: B  <= w8_L1_N4_14;
                        4: B  <= w8_L1_N5_14;
                        5: B  <= w8_L1_N6_14;
                        6: B  <= w8_L1_N7_14;
                        7: B  <= w8_L1_N8_14;
                        8: B  <= w8_L1_N9_14;
                        9: B  <= w8_L1_N10_14;
                       10: B  <= w8_L1_N11_14;
                       11: B  <= w8_L1_N12_14;
                       12: B  <= w8_L1_N13_14;
                       13: B  <= w8_L1_N14_14;
                       14: B  <= w8_L1_N15_14;
                       15: B  <= w8_L1_N16_14;
                       16: B  <= w8_L1_N17_14;
                       17: B  <= w8_L1_N18_14;
                       18: B  <= w8_L1_N19_14;
                       19: B  <= w8_L1_N20_14;
                       20: B  <= w8_L1_N21_14;
                       21: B  <= w8_L1_N22_14;
                       22: B  <= w8_L1_N23_14;
                       23: B  <= w8_L1_N24_14;
                       24: B  <= w8_L1_N25_14;
                       25: B  <= w8_L1_N26_14;
                       26: B  <= w8_L1_N27_14;
                       27: B  <= w8_L1_N28_14;
                       28: B  <= w8_L1_N29_14;
                       29: B  <= w8_L1_N30_14;
                       30: B  <= w8_L1_N31_14;
                       31: B  <= w8_L1_N32_14;
                       32: B  <= w8_L1_N33_14;
                       33: B  <= w8_L1_N34_14;
                       34: B  <= w8_L1_N35_14;
                       35: B  <= w8_L1_N36_14;
                       36: B  <= w8_L1_N37_14;
                       37: B  <= w8_L1_N38_14;
                       38: B  <= w8_L1_N39_14;
                       39: B  <= w8_L1_N40_14;
                       40: B  <= w8_L1_N41_14;
                       41: B  <= w8_L1_N42_14;
                       42: B  <= w8_L1_N43_14;
                       43: B  <= w8_L1_N44_14;
                       44: B  <= w8_L1_N45_14;
                       45: B  <= w8_L1_N46_14;
                       46: B  <= w8_L1_N47_14;
                       47: B  <= w8_L1_N48_14;
                       48: B  <= w8_L1_N49_14;
                       49: B  <= w8_L1_N50_14;
                       50: B  <= w8_L1_N51_14;
                       51: B  <= w8_L1_N52_14;
                       52: B  <= w8_L1_N53_14;
                       53: B  <= w8_L1_N54_14;
                       54: B  <= w8_L1_N55_14;
                       55: B  <= w8_L1_N56_14;
                       56: B  <= w8_L1_N57_14;
                       57: B  <= w8_L1_N58_14;
                       58: B  <= w8_L1_N59_14;
                       59: B  <= w8_L1_N60_14;
                    endcase
                end
                15: begin
                    A  <= LBP_14_fix;  //LBP_7_fix   
                    B  <= w8_L1_N1_15;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_15;
                        1: B  <= w8_L1_N2_15;
                        2: B  <= w8_L1_N3_15;
                        3: B  <= w8_L1_N4_15;
                        4: B  <= w8_L1_N5_15;
                        5: B  <= w8_L1_N6_15;
                        6: B  <= w8_L1_N7_15;
                        7: B  <= w8_L1_N8_15;
                        8: B  <= w8_L1_N9_15;
                        9: B  <= w8_L1_N10_15;
                       10: B  <= w8_L1_N11_15;
                       11: B  <= w8_L1_N12_15;
                       12: B  <= w8_L1_N13_15;
                       13: B  <= w8_L1_N14_15;
                       14: B  <= w8_L1_N15_15;
                       15: B  <= w8_L1_N16_15;
                       16: B  <= w8_L1_N17_15;
                       17: B  <= w8_L1_N18_15;
                       18: B  <= w8_L1_N19_15;
                       19: B  <= w8_L1_N20_15;
                       20: B  <= w8_L1_N21_15;
                       21: B  <= w8_L1_N22_15;
                       22: B  <= w8_L1_N23_15;
                       23: B  <= w8_L1_N24_15;
                       24: B  <= w8_L1_N25_15;
                       25: B  <= w8_L1_N26_15;
                       26: B  <= w8_L1_N27_15;
                       27: B  <= w8_L1_N28_15;
                       28: B  <= w8_L1_N29_15;
                       29: B  <= w8_L1_N30_15;
                       30: B  <= w8_L1_N31_15;
                       31: B  <= w8_L1_N32_15;
                       32: B  <= w8_L1_N33_15;
                       33: B  <= w8_L1_N34_15;
                       34: B  <= w8_L1_N35_15;
                       35: B  <= w8_L1_N36_15;
                       36: B  <= w8_L1_N37_15;
                       37: B  <= w8_L1_N38_15;
                       38: B  <= w8_L1_N39_15;
                       39: B  <= w8_L1_N40_15;
                       40: B  <= w8_L1_N41_15;
                       41: B  <= w8_L1_N42_15;
                       42: B  <= w8_L1_N43_15;
                       43: B  <= w8_L1_N44_15;
                       44: B  <= w8_L1_N45_15;
                       45: B  <= w8_L1_N46_15;
                       46: B  <= w8_L1_N47_15;
                       47: B  <= w8_L1_N48_15;
                       48: B  <= w8_L1_N49_15;
                       49: B  <= w8_L1_N50_15;
                       50: B  <= w8_L1_N51_15;
                       51: B  <= w8_L1_N52_15;
                       52: B  <= w8_L1_N53_15;
                       53: B  <= w8_L1_N54_15;
                       54: B  <= w8_L1_N55_15;
                       55: B  <= w8_L1_N56_15;
                       56: B  <= w8_L1_N57_15;
                       57: B  <= w8_L1_N58_15;
                       58: B  <= w8_L1_N59_15;
                       59: B  <= w8_L1_N60_15;
                    endcase
                end
            16: begin
                    A  <= LBP_7_fix;  //LBP_7_fix   
                    B  <= w8_L1_N1_16;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L1_N1_16;
                        1: B  <= w8_L1_N2_16;
                        2: B  <= w8_L1_N3_16;
                        3: B  <= w8_L1_N4_16;
                        4: B  <= w8_L1_N5_16;
                        5: B  <= w8_L1_N6_16;
                        6: B  <= w8_L1_N7_16;
                        7: B  <= w8_L1_N8_16;
                        8: B  <= w8_L1_N9_16;
                        9: B  <= w8_L1_N10_16;
                       10: B  <= w8_L1_N11_16;
                       11: B  <= w8_L1_N12_16;
                       12: B  <= w8_L1_N13_16;
                       13: B  <= w8_L1_N14_16;
                       14: B  <= w8_L1_N15_16;
                       15: B  <= w8_L1_N16_16;
                       16: B  <= w8_L1_N17_16;
                       17: B  <= w8_L1_N18_16;
                       18: B  <= w8_L1_N19_16;
                       19: B  <= w8_L1_N20_16;
                       20: B  <= w8_L1_N21_16;
                       21: B  <= w8_L1_N22_16;
                       22: B  <= w8_L1_N23_16;
                       23: B  <= w8_L1_N24_16;
                       24: B  <= w8_L1_N25_16;
                       25: B  <= w8_L1_N26_16;
                       26: B  <= w8_L1_N27_16;
                       27: B  <= w8_L1_N28_16;
                       28: B  <= w8_L1_N29_16;
                       29: B  <= w8_L1_N30_16;
                       30: B  <= w8_L1_N31_16;
                       31: B  <= w8_L1_N32_16;
                       32: B  <= w8_L1_N33_16;
                       33: B  <= w8_L1_N34_16;
                       34: B  <= w8_L1_N35_16;
                       35: B  <= w8_L1_N36_16;
                       36: B  <= w8_L1_N37_16;
                       37: B  <= w8_L1_N38_16;
                       38: B  <= w8_L1_N39_16;
                       39: B  <= w8_L1_N40_16;
                       40: B  <= w8_L1_N41_16;
                       41: B  <= w8_L1_N42_16;
                       42: B  <= w8_L1_N43_16;
                       43: B  <= w8_L1_N44_16;
                       44: B  <= w8_L1_N45_16;
                       45: B  <= w8_L1_N46_16;
                       46: B  <= w8_L1_N47_16;
                       47: B  <= w8_L1_N48_16;
                       48: B  <= w8_L1_N49_16;
                       49: B  <= w8_L1_N50_16;
                       50: B  <= w8_L1_N51_16;
                       51: B  <= w8_L1_N52_16;
                       52: B  <= w8_L1_N53_16;
                       53: B  <= w8_L1_N54_16;
                       54: B  <= w8_L1_N55_16;
                       55: B  <= w8_L1_N56_16;
                       56: B  <= w8_L1_N57_16;
                       57: B  <= w8_L1_N58_16;
                       58: B  <= w8_L1_N59_16;
                       59: B  <= w8_L1_N60_16;
                    endcase
                end
            endcase
            CE       <= 1;
            count    <= 0;
            nn_state <= waiting_L1_NN;
        end
        waiting_L1_NN: begin
            CE <= 1;
            if(count == 10) begin  //wait done MAC done
                NN_aggre <= P;
                if(count_input == 16)
                    nn_state    <= comp_L1_NN;
                else begin
                    count_input <= count_input + 1; //compute for next input
                    nn_state    <= start_L1_NN;
                end
            end
            else begin
               count    <= count + 1; //wait for MAC operation
               nn_state <= waiting_L1_NN;
            end
        end
        comp_L1_NN: begin
            nn_state    <= next_L1_NN;
            if(NN_aggre[58] == 1)
                NN_aggre <=59'd0;
        end
        
        next_L1_NN: begin
            if(count_NN == 59) begin
                nn_state    <= done_L1_NN;
                count_input <= 0;
                NN_aggre    <= 0;
                count       <= 0; 
            end  
            else begin
                nn_state    <= start_L1_NN;
                count_NN    <= count_NN + 1;
                count_input <= 0;
                NN_aggre    <= 0;
                count       <= 0;    
            end
            case(count_NN)
                0:  N1_L1  <= NN_aggre[48:19]; //61 --> 21.40    //31 -->  11.20  [50:20]
                1:  N2_L1  <= NN_aggre[48:19]; //50 --> 20.30    //26 -->  11.15  [40:15]
                2:  N3_L1  <= NN_aggre[48:19]; //57 --> 21.36    //29 -->  11.18  [46:18]
                3:  N4_L1  <= NN_aggre[48:19]; //59 --> 21.38    //30 -->  11.19  [48:19]
                4:  N5_L1  <= NN_aggre[48:19];
                5:  N6_L1  <= NN_aggre[48:19];
                6:  N7_L1  <= NN_aggre[48:19];
                7:  N8_L1  <= NN_aggre[48:19];
                8:  N9_L1  <= NN_aggre[48:19];
                9:  N10_L1 <= NN_aggre[48:19];
                10: N11_L1 <= NN_aggre[48:19];
                11: N12_L1 <= NN_aggre[48:19];
                12: N13_L1 <= NN_aggre[48:19];
                13: N14_L1 <= NN_aggre[48:19];
                14: N15_L1 <= NN_aggre[48:19];
                15: N16_L1 <= NN_aggre[48:19];
                16: N17_L1 <= NN_aggre[48:19];
                17: N18_L1 <= NN_aggre[48:19];
                18: N19_L1 <= NN_aggre[48:19];
                19: N20_L1 <= NN_aggre[48:19];
                20: N21_L1 <= NN_aggre[48:19];
                21: N22_L1 <= NN_aggre[48:19];
                22: N23_L1 <= NN_aggre[48:19];
                23: N24_L1 <= NN_aggre[48:19];
                24: N25_L1 <= NN_aggre[48:19];
                25: N26_L1 <= NN_aggre[48:19];
                26: N27_L1 <= NN_aggre[48:19];
                27: N28_L1 <= NN_aggre[48:19];
                28: N29_L1 <= NN_aggre[48:19];
                29: N30_L1 <= NN_aggre[48:19];
                30: N31_L1  <= NN_aggre[48:19]; //61 --> 21.40    //31 -->  11.20  [50:20]
                31: N32_L1  <= NN_aggre[48:19]; //50 --> 20.30    //26 -->  11.15  [40:15]
                32: N33_L1  <= NN_aggre[48:19]; //57 --> 21.36    //29 -->  11.18  [46:18]
                33: N34_L1  <= NN_aggre[48:19]; //59 --> 21.38    //30 -->  11.19  [48:19]
                34: N35_L1  <= NN_aggre[48:19];
                35: N36_L1  <= NN_aggre[48:19];
                36: N37_L1  <= NN_aggre[48:19];
                37: N38_L1  <= NN_aggre[48:19];
                38: N39_L1  <= NN_aggre[48:19];
                39: N40_L1 <= NN_aggre[48:19];
                40: N41_L1 <= NN_aggre[48:19];
                41: N42_L1 <= NN_aggre[48:19];
                42: N43_L1 <= NN_aggre[48:19];
                43: N44_L1 <= NN_aggre[48:19];
                44: N45_L1 <= NN_aggre[48:19];
                45: N46_L1 <= NN_aggre[48:19];
                46: N47_L1 <= NN_aggre[48:19];
                47: N48_L1 <= NN_aggre[48:19];
                48: N49_L1 <= NN_aggre[48:19];
                49: N50_L1 <= NN_aggre[48:19];
                50: N51_L1 <= NN_aggre[48:19];
                51: N52_L1 <= NN_aggre[48:19];
                52: N53_L1 <= NN_aggre[48:19];
                53: N54_L1 <= NN_aggre[48:19];
                54: N55_L1 <= NN_aggre[48:19];
                55: N56_L1 <= NN_aggre[48:19];
                56: N57_L1 <= NN_aggre[48:19];
                57: N58_L1 <= NN_aggre[48:19];
                58: N59_L1 <= NN_aggre[48:19];
                59: N60_L1 <= NN_aggre[48:19];
            endcase
        end
        done_L1_NN: begin
            nn_state    <= start_L2_NN;
            count_NN    <= 0;
        end

       start_L2_NN: begin
            case(count_input)
                0: begin
                    A  <= N1_L1;
                    case(count_NN)
                        0: begin B  <= w8_L2_N1_0;   C  <= b_L2_N1; end
                        1: begin B  <= w8_L2_N2_0;   C  <= b_L2_N2; end
                        2: begin B  <= w8_L2_N3_0;   C  <= b_L2_N3; end
                        3: begin B  <= w8_L2_N4_0;   C  <= b_L2_N4; end
                        4: begin B  <= w8_L2_N5_0;   C  <= b_L2_N5; end
                        5: begin B  <= w8_L2_N6_0;   C  <= b_L2_N6; end
                        6: begin B  <= w8_L2_N7_0;   C  <= b_L2_N7; end
                        7: begin B  <= w8_L2_N8_0;   C  <= b_L2_N8; end
                        8: begin B  <= w8_L2_N9_0;   C  <= b_L2_N9; end
                        9: begin B  <= w8_L2_N10_0;  C  <= b_L2_N10; end
                        10:begin B  <= w8_L2_N11_0;  C  <= b_L2_N11; end
                        11:begin B  <= w8_L2_N12_0;  C  <= b_L2_N12; end
                        12:begin B  <= w8_L2_N13_0;  C  <= b_L2_N13; end
                        13:begin B  <= w8_L2_N14_0;  C  <= b_L2_N14; end
                        14:begin B  <= w8_L2_N15_0;  C  <= b_L2_N15; end
                        15:begin B  <= w8_L2_N16_0;  C  <= b_L2_N16; end
                        16:begin B  <= w8_L2_N17_0;  C  <= b_L2_N17; end
                        17:begin B  <= w8_L2_N18_0;  C  <= b_L2_N18; end
                        18:begin B  <= w8_L2_N19_0;  C  <= b_L2_N19; end
                        19:begin B  <= w8_L2_N20_0;  C  <= b_L2_N20; end
                    endcase
                end
                1: begin
                    A  <= N2_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_1;
                        1: B  <= w8_L2_N2_1;
                        2: B  <= w8_L2_N3_1;
                        3: B  <= w8_L2_N4_1;
                        4: B  <= w8_L2_N5_1;
                        5: B  <= w8_L2_N6_1;
                        6: B  <= w8_L2_N7_1;
                        7: B  <= w8_L2_N8_1;
                        8: B  <= w8_L2_N9_1;
                        9: B  <= w8_L2_N10_1;
                        10:B  <= w8_L2_N11_1;
                        11:B  <= w8_L2_N12_1;
                        12:B  <= w8_L2_N13_1;
                        13:B  <= w8_L2_N14_1;
                        14:B  <= w8_L2_N15_1;
                        15:B  <= w8_L2_N16_1;
                        16:B  <= w8_L2_N17_1;
                        17:B  <= w8_L2_N18_1;
                        18:B  <= w8_L2_N19_1;
                        19:B  <= w8_L2_N20_1;
                    endcase
                end
                2: begin
                    A  <= N3_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_2;
                        1: B  <= w8_L2_N2_2;
                        2: B  <= w8_L2_N3_2;
                        3: B  <= w8_L2_N4_2;
                        4: B  <= w8_L2_N5_2;
                        5: B  <= w8_L2_N6_2;
                        6: B  <= w8_L2_N7_2;
                        7: B  <= w8_L2_N8_2;
                        8: B  <= w8_L2_N9_2; 
                        9: B  <= w8_L2_N10_2;
                        10:B  <= w8_L2_N11_2;
                        11:B  <= w8_L2_N12_2;
                        12:B  <= w8_L2_N13_2;
                        13:B  <= w8_L2_N14_2;
                        14:B  <= w8_L2_N15_2;
                        15:B  <= w8_L2_N16_2;
                        16:B  <= w8_L2_N17_2;
                        17:B  <= w8_L2_N18_2;
                        18:B  <= w8_L2_N19_2;
                        19:B  <= w8_L2_N20_2;
                    endcase
                end
                3: begin
                    A  <= N4_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_3;
                        1: B  <= w8_L2_N2_3;
                        2: B  <= w8_L2_N3_3;
                        3: B  <= w8_L2_N4_3;
                        4: B  <= w8_L2_N5_3;
                        5: B  <= w8_L2_N6_3;
                        6: B  <= w8_L2_N7_3;
                        7: B  <= w8_L2_N8_3;
                        8: B  <= w8_L2_N9_3;
                        9: B  <= w8_L2_N10_3;
                        10:B  <= w8_L2_N11_3;
                        11:B  <= w8_L2_N12_3;
                        12:B  <= w8_L2_N13_3;
                        13:B  <= w8_L2_N14_3;
                        14:B  <= w8_L2_N15_3;
                        15:B  <= w8_L2_N16_3;
                        16:B  <= w8_L2_N17_3;
                        17:B  <= w8_L2_N18_3;
                        18:B  <= w8_L2_N19_3;
                        19:B  <= w8_L2_N20_3;
                    endcase
                end
                4: begin
                    A  <= N5_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_4;
                        1: B  <= w8_L2_N2_4;
                        2: B  <= w8_L2_N3_4;
                        3: B  <= w8_L2_N4_4;
                        4: B  <= w8_L2_N5_4;
                        5: B  <= w8_L2_N6_4;
                        6: B  <= w8_L2_N7_4;
                        7: B  <= w8_L2_N8_4;
                        8: B  <= w8_L2_N9_4;
                        9: B  <= w8_L2_N10_4;
                        10:B  <= w8_L2_N11_4;
                        11:B  <= w8_L2_N12_4;
                        12:B  <= w8_L2_N13_4;
                        13:B  <= w8_L2_N14_4;
                        14:B  <= w8_L2_N15_4;
                        15:B  <= w8_L2_N16_4;
                        16:B  <= w8_L2_N17_4;
                        17:B  <= w8_L2_N18_4;
                        18:B  <= w8_L2_N19_4;
                        19:B  <= w8_L2_N20_4;
                    endcase
                end
                5: begin
                    A  <= N6_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_5;
                        1: B  <= w8_L2_N2_5;
                        2: B  <= w8_L2_N3_5;
                        3: B  <= w8_L2_N4_5;
                        4: B  <= w8_L2_N5_5;
                        5: B  <= w8_L2_N6_5;
                        6: B  <= w8_L2_N7_5;
                        7: B  <= w8_L2_N8_5;
                        8: B  <= w8_L2_N9_5;
                        9: B  <= w8_L2_N10_5;
                        10:B  <= w8_L2_N11_5;
                        11:B  <= w8_L2_N12_5;
                        12:B  <= w8_L2_N13_5;
                        13:B  <= w8_L2_N14_5;
                        14:B  <= w8_L2_N15_5;
                        15:B  <= w8_L2_N16_5;
                        16:B  <= w8_L2_N17_5;
                        17:B  <= w8_L2_N18_5;
                        18:B  <= w8_L2_N19_5;
                        19:B  <= w8_L2_N20_5;
                    endcase
                end
                6: begin
                    A  <= N7_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_6;
                        1: B  <= w8_L2_N2_6;
                        2: B  <= w8_L2_N3_6;
                        3: B  <= w8_L2_N4_6;
                        4: B  <= w8_L2_N5_6;
                        5: B  <= w8_L2_N6_6;
                        6: B  <= w8_L2_N7_6;
                        7: B  <= w8_L2_N8_6;
                        8: B  <= w8_L2_N9_6;
                        9: B  <= w8_L2_N10_6;
                        10:B  <= w8_L2_N11_6;
                        11:B  <= w8_L2_N12_6;
                        12:B  <= w8_L2_N13_6;
                        13:B  <= w8_L2_N14_6;
                        14:B  <= w8_L2_N15_6;
                        15:B  <= w8_L2_N16_6;
                        16:B  <= w8_L2_N17_6;
                        17:B  <= w8_L2_N18_6;
                        18:B  <= w8_L2_N19_6;
                        19:B  <= w8_L2_N20_6;
                    endcase
                end
                7: begin
                    A  <= N8_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_7;
                        1: B  <= w8_L2_N2_7;
                        2: B  <= w8_L2_N3_7;
                        3: B  <= w8_L2_N4_7;
                        4: B  <= w8_L2_N5_7;
                        5: B  <= w8_L2_N6_7;
                        6: B  <= w8_L2_N7_7;
                        7: B  <= w8_L2_N8_7;
                        8: B  <= w8_L2_N9_7;
                        9: B  <= w8_L2_N10_7;
                        10:B  <= w8_L2_N11_7;
                        11:B  <= w8_L2_N12_7;
                        12:B  <= w8_L2_N13_7;
                        13:B  <= w8_L2_N14_7;
                        14:B  <= w8_L2_N15_7;
                        15:B  <= w8_L2_N16_7;
                        16:B  <= w8_L2_N17_7;
                        17:B  <= w8_L2_N18_7;
                        18:B  <= w8_L2_N19_7;
                        19:B  <= w8_L2_N20_7;
                    endcase
                end
                8: begin
                    A  <= N9_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_8;
                        1: B  <= w8_L2_N2_8;
                        2: B  <= w8_L2_N3_8;
                        3: B  <= w8_L2_N4_8;
                        4: B  <= w8_L2_N5_8;
                        5: B  <= w8_L2_N6_8;
                        6: B  <= w8_L2_N7_8;
                        7: B  <= w8_L2_N8_8;
                        8: B  <= w8_L2_N9_8;
                        9: B  <= w8_L2_N10_8;
                        10:B  <= w8_L2_N11_8;
                        11:B  <= w8_L2_N12_8;
                        12:B  <= w8_L2_N13_8;
                        13:B  <= w8_L2_N14_8;
                        14:B  <= w8_L2_N15_8;
                        15:B  <= w8_L2_N16_8;
                        16:B  <= w8_L2_N17_8;
                        17:B  <= w8_L2_N18_8;
                        18:B  <= w8_L2_N19_8;
                        19:B  <= w8_L2_N20_8;
                    endcase
                end
                9: begin
                    A  <= N10_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_9;
                        1: B  <= w8_L2_N2_9;
                        2: B  <= w8_L2_N3_9;
                        3: B  <= w8_L2_N4_9;
                        4: B  <= w8_L2_N5_9;
                        5: B  <= w8_L2_N6_9;
                        6: B  <= w8_L2_N7_9;
                        7: B  <= w8_L2_N8_9;
                        8: B  <= w8_L2_N9_9;
                        9: B  <= w8_L2_N10_9;
                        10:B  <= w8_L2_N11_9;
                        11:B  <= w8_L2_N12_9;
                        12:B  <= w8_L2_N13_9;
                        13:B  <= w8_L2_N14_9;
                        14:B  <= w8_L2_N15_9;
                        15:B  <= w8_L2_N16_9;
                        16:B  <= w8_L2_N17_9;
                        17:B  <= w8_L2_N18_9;
                        18:B  <= w8_L2_N19_9;
                        19:B  <= w8_L2_N20_9;
                    endcase
                end
                10: begin
                    A  <= N11_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_10;
                        1: B  <= w8_L2_N2_10;
                        2: B  <= w8_L2_N3_10;
                        3: B  <= w8_L2_N4_10;
                        4: B  <= w8_L2_N5_10;
                        5: B  <= w8_L2_N6_10;
                        6: B  <= w8_L2_N7_10;
                        7: B  <= w8_L2_N8_10;
                        8: B  <= w8_L2_N9_10;
                        9: B  <= w8_L2_N10_10;
                        10:B  <= w8_L2_N11_10;
                        11:B  <= w8_L2_N12_10;
                        12:B  <= w8_L2_N13_10;
                        13:B  <= w8_L2_N14_10;
                        14:B  <= w8_L2_N15_10;
                        15:B  <= w8_L2_N16_10;
                        16:B  <= w8_L2_N17_10;
                        17:B  <= w8_L2_N18_10;
                        18:B  <= w8_L2_N19_10;
                        19:B  <= w8_L2_N20_10;
                    endcase
                end
                11: begin
                    A  <= N12_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_11;
                        1: B  <= w8_L2_N2_11;
                        2: B  <= w8_L2_N3_11;
                        3: B  <= w8_L2_N4_11;
                        4: B  <= w8_L2_N5_11;
                        5: B  <= w8_L2_N6_11;
                        6: B  <= w8_L2_N7_11;
                        7: B  <= w8_L2_N8_11;
                        8: B  <= w8_L2_N9_11;
                        9: B  <= w8_L2_N10_11;
                        10:B  <= w8_L2_N11_11;
                        11:B  <= w8_L2_N12_11;
                        12:B  <= w8_L2_N13_11;
                        13:B  <= w8_L2_N14_11;
                        14:B  <= w8_L2_N15_11;
                        15:B  <= w8_L2_N16_11;
                        16:B  <= w8_L2_N17_11;
                        17:B  <= w8_L2_N18_11;
                        18:B  <= w8_L2_N19_11;
                        19:B  <= w8_L2_N20_11;
                    endcase
                end
                12: begin
                    A  <= N13_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_12;
                        1: B  <= w8_L2_N2_12;
                        2: B  <= w8_L2_N3_12;
                        3: B  <= w8_L2_N4_12;
                        4: B  <= w8_L2_N5_12;
                        5: B  <= w8_L2_N6_12;
                        6: B  <= w8_L2_N7_12;
                        7: B  <= w8_L2_N8_12;
                        8: B  <= w8_L2_N9_12;
                        9: B  <= w8_L2_N10_12;
                        10:B  <= w8_L2_N11_12;
                        11:B  <= w8_L2_N12_12;
                        12:B  <= w8_L2_N13_12;
                        13:B  <= w8_L2_N14_12;
                        14:B  <= w8_L2_N15_12;
                        15:B  <= w8_L2_N16_12;
                        16:B  <= w8_L2_N17_12;
                        17:B  <= w8_L2_N18_12;
                        18:B  <= w8_L2_N19_12;
                        19:B  <= w8_L2_N20_12;
                    endcase
                end
                13: begin
                    A  <= N14_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_13;
                        1: B  <= w8_L2_N2_13;
                        2: B  <= w8_L2_N3_13;
                        3: B  <= w8_L2_N4_13;
                        4: B  <= w8_L2_N5_13;
                        5: B  <= w8_L2_N6_13;
                        6: B  <= w8_L2_N7_13;
                        7: B  <= w8_L2_N8_13;
                        8: B  <= w8_L2_N9_13;
                        9: B  <= w8_L2_N10_13;
                        10:B  <= w8_L2_N11_13;
                        11:B  <= w8_L2_N12_13;
                        12:B  <= w8_L2_N13_13;
                        13:B  <= w8_L2_N14_13;
                        14:B  <= w8_L2_N15_13;
                        15:B  <= w8_L2_N16_13;
                        16:B  <= w8_L2_N17_13;
                        17:B  <= w8_L2_N18_13;
                        18:B  <= w8_L2_N19_13;
                        19:B  <= w8_L2_N20_13;
                    endcase
                end
                14: begin
                    A  <= N15_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_14;
                        1: B  <= w8_L2_N2_14;
                        2: B  <= w8_L2_N3_14;
                        3: B  <= w8_L2_N4_14;
                        4: B  <= w8_L2_N5_14;
                        5: B  <= w8_L2_N6_14;
                        6: B  <= w8_L2_N7_14;
                        7: B  <= w8_L2_N8_14;
                        8: B  <= w8_L2_N9_14;
                        9: B  <= w8_L2_N10_14;
                        10:B  <= w8_L2_N11_14;
                        11:B  <= w8_L2_N12_14;
                        12:B  <= w8_L2_N13_14;
                        13:B  <= w8_L2_N14_14;
                        14:B  <= w8_L2_N15_14;
                        15:B  <= w8_L2_N16_14;
                        16:B  <= w8_L2_N17_14;
                        17:B  <= w8_L2_N18_14;
                        18:B  <= w8_L2_N19_14;
                        19:B  <= w8_L2_N20_14;
                    endcase
                end
                15: begin
                    A  <= N16_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_15;
                        1: B  <= w8_L2_N2_15;
                        2: B  <= w8_L2_N3_15;
                        3: B  <= w8_L2_N4_15;
                        4: B  <= w8_L2_N5_15;
                        5: B  <= w8_L2_N6_15;
                        6: B  <= w8_L2_N7_15;
                        7: B  <= w8_L2_N8_15;
                        8: B  <= w8_L2_N9_15;
                        9: B  <= w8_L2_N10_15;
                        10:B  <= w8_L2_N11_15;
                        11:B  <= w8_L2_N12_15;
                        12:B  <= w8_L2_N13_15;
                        13:B  <= w8_L2_N14_15;
                        14:B  <= w8_L2_N15_15;
                        15:B  <= w8_L2_N16_15;
                        16:B  <= w8_L2_N17_15;
                        17:B  <= w8_L2_N18_15;
                        18:B  <= w8_L2_N19_15;
                        19:B  <= w8_L2_N20_15;
                    endcase
                end
                16: begin
                    A  <= N17_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_16;
                        1: B  <= w8_L2_N2_16;
                        2: B  <= w8_L2_N3_16;
                        3: B  <= w8_L2_N4_16;
                        4: B  <= w8_L2_N5_16;
                        5: B  <= w8_L2_N6_16;
                        6: B  <= w8_L2_N7_16;
                        7: B  <= w8_L2_N8_16;
                        8: B  <= w8_L2_N9_16;
                        9: B  <= w8_L2_N10_16;
                        10:B  <= w8_L2_N11_16;
                        11:B  <= w8_L2_N12_16;
                        12:B  <= w8_L2_N13_16;
                        13:B  <= w8_L2_N14_16;
                        14:B  <= w8_L2_N15_16;
                        15:B  <= w8_L2_N16_16;
                        16:B  <= w8_L2_N17_16;
                        17:B  <= w8_L2_N18_16;
                        18:B  <= w8_L2_N19_16;
                        19:B  <= w8_L2_N20_16;
                    endcase
                end
                17: begin
                    A  <= N18_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_17;
                        1: B  <= w8_L2_N2_17;
                        2: B  <= w8_L2_N3_17;
                        3: B  <= w8_L2_N4_17;
                        4: B  <= w8_L2_N5_17;
                        5: B  <= w8_L2_N6_17;
                        6: B  <= w8_L2_N7_17;
                        7: B  <= w8_L2_N8_17;
                        8: B  <= w8_L2_N9_17;
                        9: B  <= w8_L2_N10_17;
                        10:B  <= w8_L2_N11_17;
                        11:B  <= w8_L2_N12_17;
                        12:B  <= w8_L2_N13_17;
                        13:B  <= w8_L2_N14_17;
                        14:B  <= w8_L2_N15_17;
                        15:B  <= w8_L2_N16_17;
                        16:B  <= w8_L2_N17_17;
                        17:B  <= w8_L2_N18_17;
                        18:B  <= w8_L2_N19_17;
                        19:B  <= w8_L2_N20_17;
                    endcase
                end
                18: begin
                    A  <= N19_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_18;
                        1: B  <= w8_L2_N2_18;
                        2: B  <= w8_L2_N3_18;
                        3: B  <= w8_L2_N4_18;
                        4: B  <= w8_L2_N5_18;
                        5: B  <= w8_L2_N6_18;
                        6: B  <= w8_L2_N7_18;
                        7: B  <= w8_L2_N8_18;
                        8: B  <= w8_L2_N9_18;
                        9: B  <= w8_L2_N10_18;
                        10:B  <= w8_L2_N11_18;
                        11:B  <= w8_L2_N12_18;
                        12:B  <= w8_L2_N13_18;
                        13:B  <= w8_L2_N14_18;
                        14:B  <= w8_L2_N15_18;
                        15:B  <= w8_L2_N16_18;
                        16:B  <= w8_L2_N17_18;
                        17:B  <= w8_L2_N18_18;
                        18:B  <= w8_L2_N19_18;
                        19:B  <= w8_L2_N20_18;
                    endcase
                end
                19: begin
                    A  <= N20_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_19;
                        1: B  <= w8_L2_N2_19;
                        2: B  <= w8_L2_N3_19;
                        3: B  <= w8_L2_N4_19;
                        4: B  <= w8_L2_N5_19;
                        5: B  <= w8_L2_N6_19;
                        6: B  <= w8_L2_N7_19;
                        7: B  <= w8_L2_N8_19;
                        8: B  <= w8_L2_N9_19;
                        9: B  <= w8_L2_N10_19;
                        10:B  <= w8_L2_N11_19;
                        11:B  <= w8_L2_N12_19;
                        12:B  <= w8_L2_N13_19;
                        13:B  <= w8_L2_N14_19;
                        14:B  <= w8_L2_N15_19;
                        15:B  <= w8_L2_N16_19;
                        16:B  <= w8_L2_N17_19;
                        17:B  <= w8_L2_N18_19;
                        18:B  <= w8_L2_N19_19;
                        19:B  <= w8_L2_N20_19;
                    endcase
                end
                20: begin
                    A  <= N21_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_20;
                        1: B  <= w8_L2_N2_20;
                        2: B  <= w8_L2_N3_20;
                        3: B  <= w8_L2_N4_20;
                        4: B  <= w8_L2_N5_20;
                        5: B  <= w8_L2_N6_20;
                        6: B  <= w8_L2_N7_20;
                        7: B  <= w8_L2_N8_20;
                        8: B  <= w8_L2_N9_20;
                        9: B  <= w8_L2_N10_20;
                        10:B  <= w8_L2_N11_20;
                        11:B  <= w8_L2_N12_20;
                        12:B  <= w8_L2_N13_20;
                        13:B  <= w8_L2_N14_20;
                        14:B  <= w8_L2_N15_20;
                        15:B  <= w8_L2_N16_20;
                        16:B  <= w8_L2_N17_20;
                        17:B  <= w8_L2_N18_20;
                        18:B  <= w8_L2_N19_20;
                        19:B  <= w8_L2_N20_20;
                    endcase
                end
                21: begin
                    A  <= N22_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_21;
                        1: B  <= w8_L2_N2_21;
                        2: B  <= w8_L2_N3_21;
                        3: B  <= w8_L2_N4_21;
                        4: B  <= w8_L2_N5_21;
                        5: B  <= w8_L2_N6_21;
                        6: B  <= w8_L2_N7_21;
                        7: B  <= w8_L2_N8_21;
                        8: B  <= w8_L2_N9_21;
                        9: B  <= w8_L2_N10_21;
                        10:B  <= w8_L2_N11_21;
                        11:B  <= w8_L2_N12_21;
                        12:B  <= w8_L2_N13_21;
                        13:B  <= w8_L2_N14_21;
                        14:B  <= w8_L2_N15_21;
                        15:B  <= w8_L2_N16_21;
                        16:B  <= w8_L2_N17_21;
                        17:B  <= w8_L2_N18_21;
                        18:B  <= w8_L2_N19_21;
                        19:B  <= w8_L2_N20_21;
                    endcase
                end
                22: begin
                    A  <= N23_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_22;
                        1: B  <= w8_L2_N2_22;
                        2: B  <= w8_L2_N3_22;
                        3: B  <= w8_L2_N4_22;
                        4: B  <= w8_L2_N5_22;
                        5: B  <= w8_L2_N6_22;
                        6: B  <= w8_L2_N7_22;
                        7: B  <= w8_L2_N8_22;
                        8: B  <= w8_L2_N9_22;
                        9: B  <= w8_L2_N10_22;
                        10:B  <= w8_L2_N11_22;
                        11:B  <= w8_L2_N12_22;
                        12:B  <= w8_L2_N13_22;
                        13:B  <= w8_L2_N14_22;
                        14:B  <= w8_L2_N15_22;
                        15:B  <= w8_L2_N16_22;
                        16:B  <= w8_L2_N17_22;
                        17:B  <= w8_L2_N18_22;
                        18:B  <= w8_L2_N19_22;
                        19:B  <= w8_L2_N20_22;
                    endcase
                end
                23: begin
                    A  <= N24_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_23;
                        1: B  <= w8_L2_N2_23;
                        2: B  <= w8_L2_N3_23;
                        3: B  <= w8_L2_N4_23;
                        4: B  <= w8_L2_N5_23;
                        5: B  <= w8_L2_N6_23;
                        6: B  <= w8_L2_N7_23;
                        7: B  <= w8_L2_N8_23;
                        8: B  <= w8_L2_N9_23;
                        9: B  <= w8_L2_N10_23;
                        10:B  <= w8_L2_N11_23;
                        11:B  <= w8_L2_N12_23;
                        12:B  <= w8_L2_N13_23;
                        13:B  <= w8_L2_N14_23;
                        14:B  <= w8_L2_N15_23;
                        15:B  <= w8_L2_N16_23;
                        16:B  <= w8_L2_N17_23;
                        17:B  <= w8_L2_N18_23;
                        18:B  <= w8_L2_N19_23;
                        19:B  <= w8_L2_N20_23;
                    endcase
                end
                24: begin
                    A  <= N25_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_24;
                        1: B  <= w8_L2_N2_24;
                        2: B  <= w8_L2_N3_24;
                        3: B  <= w8_L2_N4_24;
                        4: B  <= w8_L2_N5_24;
                        5: B  <= w8_L2_N6_24;
                        6: B  <= w8_L2_N7_24;
                        7: B  <= w8_L2_N8_24;
                        8: B  <= w8_L2_N9_24;
                        9: B  <= w8_L2_N10_24;
                        10:B  <= w8_L2_N11_24;
                        11:B  <= w8_L2_N12_24;
                        12:B  <= w8_L2_N13_24;
                        13:B  <= w8_L2_N14_24;
                        14:B  <= w8_L2_N15_24;
                        15:B  <= w8_L2_N16_24;
                        16:B  <= w8_L2_N17_24;
                        17:B  <= w8_L2_N18_24;
                        18:B  <= w8_L2_N19_24;
                        19:B  <= w8_L2_N20_24;
                    endcase
                end
                25: begin
                    A  <= N26_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_25;
                        1: B  <= w8_L2_N2_25;
                        2: B  <= w8_L2_N3_25;
                        3: B  <= w8_L2_N4_25;
                        4: B  <= w8_L2_N5_25;
                        5: B  <= w8_L2_N6_25;
                        6: B  <= w8_L2_N7_25;
                        7: B  <= w8_L2_N8_25;
                        8: B  <= w8_L2_N9_25;
                        9: B  <= w8_L2_N10_25;
                        10:B  <= w8_L2_N11_25;
                        11:B  <= w8_L2_N12_25;
                        12:B  <= w8_L2_N13_25;
                        13:B  <= w8_L2_N14_25;
                        14:B  <= w8_L2_N15_25;
                        15:B  <= w8_L2_N16_25;
                        16:B  <= w8_L2_N17_25;
                        17:B  <= w8_L2_N18_25;
                        18:B  <= w8_L2_N19_25;
                        19:B  <= w8_L2_N20_25;
                    endcase
                end
                26: begin
                    A  <= N27_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_26;
                        1: B  <= w8_L2_N2_26;
                        2: B  <= w8_L2_N3_26;
                        3: B  <= w8_L2_N4_26;
                        4: B  <= w8_L2_N5_26;
                        5: B  <= w8_L2_N6_26;
                        6: B  <= w8_L2_N7_26;
                        7: B  <= w8_L2_N8_26;
                        8: B  <= w8_L2_N9_26;
                        9: B  <= w8_L2_N10_26;
                        10:B  <= w8_L2_N11_26;
                        11:B  <= w8_L2_N12_26;
                        12:B  <= w8_L2_N13_26;
                        13:B  <= w8_L2_N14_26;
                        14:B  <= w8_L2_N15_26;
                        15:B  <= w8_L2_N16_26;
                        16:B  <= w8_L2_N17_26;
                        17:B  <= w8_L2_N18_26;
                        18:B  <= w8_L2_N19_26;
                        19:B  <= w8_L2_N20_26;
                    endcase
                end
                27: begin
                    A  <= N28_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_27;
                        1: B  <= w8_L2_N2_27;
                        2: B  <= w8_L2_N3_27;
                        3: B  <= w8_L2_N4_27;
                        4: B  <= w8_L2_N5_27;
                        5: B  <= w8_L2_N6_27;
                        6: B  <= w8_L2_N7_27;
                        7: B  <= w8_L2_N8_27;
                        8: B  <= w8_L2_N9_27;
                        9: B  <= w8_L2_N10_27;
                        10:B  <= w8_L2_N11_27;
                        11:B  <= w8_L2_N12_27;
                        12:B  <= w8_L2_N13_27;
                        13:B  <= w8_L2_N14_27;
                        14:B  <= w8_L2_N15_27;
                        15:B  <= w8_L2_N16_27;
                        16:B  <= w8_L2_N17_27;
                        17:B  <= w8_L2_N18_27;
                        18:B  <= w8_L2_N19_27;
                        19:B  <= w8_L2_N20_27;
                    endcase
                end
                28: begin
                    A  <= N29_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_28;
                        1: B  <= w8_L2_N2_28;
                        2: B  <= w8_L2_N3_28;
                        3: B  <= w8_L2_N4_28;
                        4: B  <= w8_L2_N5_28;
                        5: B  <= w8_L2_N6_28;
                        6: B  <= w8_L2_N7_28;
                        7: B  <= w8_L2_N8_28;
                        8: B  <= w8_L2_N9_28;
                        9: B  <= w8_L2_N10_28;
                        10:B  <= w8_L2_N11_28;
                        11:B  <= w8_L2_N12_28;
                        12:B  <= w8_L2_N13_28;
                        13:B  <= w8_L2_N14_28;
                        14:B  <= w8_L2_N15_28;
                        15:B  <= w8_L2_N16_28;
                        16:B  <= w8_L2_N17_28;
                        17:B  <= w8_L2_N18_28;
                        18:B  <= w8_L2_N19_28;
                        19:B  <= w8_L2_N20_28;
                    endcase
                end
                29: begin
                    A  <= N30_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <= w8_L2_N1_29;
                        1: B  <= w8_L2_N2_29;
                        2: B  <= w8_L2_N3_29;
                        3: B  <= w8_L2_N4_29;
                        4: B  <= w8_L2_N5_29;
                        5: B  <= w8_L2_N6_29;
                        6: B  <= w8_L2_N7_29;
                        7: B  <= w8_L2_N8_29;
                        8: B  <= w8_L2_N9_29;
                        9: B  <= w8_L2_N10_29;
                        10:B  <= w8_L2_N11_29;
                        11:B  <= w8_L2_N12_29;
                        12:B  <= w8_L2_N13_29;
                        13:B  <= w8_L2_N14_29;
                        14:B  <= w8_L2_N15_29;
                        15:B  <= w8_L2_N16_29;
                        16:B  <= w8_L2_N17_29;
                        17:B  <= w8_L2_N18_29;
                        18:B  <= w8_L2_N19_29;
                        19:B  <= w8_L2_N20_29;
                    endcase
                end
                30: begin
                    A  <= N31_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_30;
                        1: B  <=  w8_L2_N2_30;
                        2: B  <=  w8_L2_N3_30;
                        3: B  <=  w8_L2_N4_30;
                        4: B  <=  w8_L2_N5_30;
                        5: B  <=  w8_L2_N6_30;
                        6: B  <=  w8_L2_N7_30;
                        7: B  <=  w8_L2_N8_30;
                        8: B  <=  w8_L2_N9_30;
                        9: B  <= w8_L2_N10_30;
                        10:B  <= w8_L2_N11_30;
                        11:B  <= w8_L2_N12_30;
                        12:B  <= w8_L2_N13_30;
                        13:B  <= w8_L2_N14_30;
                        14:B  <= w8_L2_N15_30;
                        15:B  <= w8_L2_N16_30;
                        16:B  <= w8_L2_N17_30;
                        17:B  <= w8_L2_N18_30;
                        18:B  <= w8_L2_N19_30;
                        19:B  <= w8_L2_N20_30;
                    endcase
                end
               31: begin
                    A  <= N32_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_31;
                        1: B  <=  w8_L2_N2_31;
                        2: B  <=  w8_L2_N3_31;
                        3: B  <=  w8_L2_N4_31;
                        4: B  <=  w8_L2_N5_31;
                        5: B  <=  w8_L2_N6_31;
                        6: B  <=  w8_L2_N7_31;
                        7: B  <=  w8_L2_N8_31;
                        8: B  <=  w8_L2_N9_31;
                        9: B  <= w8_L2_N10_31;
                        10:B  <= w8_L2_N11_31;
                        11:B  <= w8_L2_N12_31;
                        12:B  <= w8_L2_N13_31;
                        13:B  <= w8_L2_N14_31;
                        14:B  <= w8_L2_N15_31;
                        15:B  <= w8_L2_N16_31;
                        16:B  <= w8_L2_N17_31;
                        17:B  <= w8_L2_N18_31;
                        18:B  <= w8_L2_N19_31;
                        19:B  <= w8_L2_N20_31;
                    endcase
                end

               32: begin
                    A  <= N33_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_32;
                        1: B  <=  w8_L2_N2_32;
                        2: B  <=  w8_L2_N3_32;
                        3: B  <=  w8_L2_N4_32;
                        4: B  <=  w8_L2_N5_32;
                        5: B  <=  w8_L2_N6_32;
                        6: B  <=  w8_L2_N7_32;
                        7: B  <=  w8_L2_N8_32;
                        8: B  <=  w8_L2_N9_32;
                        9: B  <= w8_L2_N10_32;
                        10:B  <= w8_L2_N11_32;
                        11:B  <= w8_L2_N12_32;
                        12:B  <= w8_L2_N13_32;
                        13:B  <= w8_L2_N14_32;
                        14:B  <= w8_L2_N15_32;
                        15:B  <= w8_L2_N16_32;
                        16:B  <= w8_L2_N17_32;
                        17:B  <= w8_L2_N18_32;
                        18:B  <= w8_L2_N19_32;
                        19:B  <= w8_L2_N20_32;
                    endcase
                end

               33: begin
                    A  <= N34_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_33;
                        1: B  <=  w8_L2_N2_33;
                        2: B  <=  w8_L2_N3_33;
                        3: B  <=  w8_L2_N4_33;
                        4: B  <=  w8_L2_N5_33;
                        5: B  <=  w8_L2_N6_33;
                        6: B  <=  w8_L2_N7_33;
                        7: B  <=  w8_L2_N8_33;
                        8: B  <=  w8_L2_N9_33;
                        9: B  <= w8_L2_N10_33;
                        10:B  <= w8_L2_N11_33;
                        11:B  <= w8_L2_N12_33;
                        12:B  <= w8_L2_N13_33;
                        13:B  <= w8_L2_N14_33;
                        14:B  <= w8_L2_N15_33;
                        15:B  <= w8_L2_N16_33;
                        16:B  <= w8_L2_N17_33;
                        17:B  <= w8_L2_N18_33;
                        18:B  <= w8_L2_N19_33;
                        19:B  <= w8_L2_N20_33;
                    endcase
                end

               34: begin
                    A  <= N35_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_34;
                        1: B  <=  w8_L2_N2_34;
                        2: B  <=  w8_L2_N3_34;
                        3: B  <=  w8_L2_N4_34;
                        4: B  <=  w8_L2_N5_34;
                        5: B  <=  w8_L2_N6_34;
                        6: B  <=  w8_L2_N7_34;
                        7: B  <=  w8_L2_N8_34;
                        8: B  <=  w8_L2_N9_34;
                        9: B  <= w8_L2_N10_34;
                        10:B  <= w8_L2_N11_34;
                        11:B  <= w8_L2_N12_34;
                        12:B  <= w8_L2_N13_34;
                        13:B  <= w8_L2_N14_34;
                        14:B  <= w8_L2_N15_34;
                        15:B  <= w8_L2_N16_34;
                        16:B  <= w8_L2_N17_34;
                        17:B  <= w8_L2_N18_34;
                        18:B  <= w8_L2_N19_34;
                        19:B  <= w8_L2_N20_34;
                    endcase
                end

               35: begin
                    A  <= N36_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_35;
                        1: B  <=  w8_L2_N2_35;
                        2: B  <=  w8_L2_N3_35;
                        3: B  <=  w8_L2_N4_35;
                        4: B  <=  w8_L2_N5_35;
                        5: B  <=  w8_L2_N6_35;
                        6: B  <=  w8_L2_N7_35;
                        7: B  <=  w8_L2_N8_35;
                        8: B  <=  w8_L2_N9_35;
                        9: B  <= w8_L2_N10_35;
                        10:B  <= w8_L2_N11_35;
                        11:B  <= w8_L2_N12_35;
                        12:B  <= w8_L2_N13_35;
                        13:B  <= w8_L2_N14_35;
                        14:B  <= w8_L2_N15_35;
                        15:B  <= w8_L2_N16_35;
                        16:B  <= w8_L2_N17_35;
                        17:B  <= w8_L2_N18_35;
                        18:B  <= w8_L2_N19_35;
                        19:B  <= w8_L2_N20_35;
                    endcase
                end

               36: begin
                    A  <= N37_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_36;
                        1: B  <=  w8_L2_N2_36;
                        2: B  <=  w8_L2_N3_36;
                        3: B  <=  w8_L2_N4_36;
                        4: B  <=  w8_L2_N5_36;
                        5: B  <=  w8_L2_N6_36;
                        6: B  <=  w8_L2_N7_36;
                        7: B  <=  w8_L2_N8_36;
                        8: B  <=  w8_L2_N9_36;
                        9: B  <= w8_L2_N10_36;
                        10:B  <= w8_L2_N11_36;
                        11:B  <= w8_L2_N12_36;
                        12:B  <= w8_L2_N13_36;
                        13:B  <= w8_L2_N14_36;
                        14:B  <= w8_L2_N15_36;
                        15:B  <= w8_L2_N16_36;
                        16:B  <= w8_L2_N17_36;
                        17:B  <= w8_L2_N18_36;
                        18:B  <= w8_L2_N19_36;
                        19:B  <= w8_L2_N20_36;
                    endcase
                end

               37: begin
                    A  <= N38_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_37;
                        1: B  <=  w8_L2_N2_37;
                        2: B  <=  w8_L2_N3_37;
                        3: B  <=  w8_L2_N4_37;
                        4: B  <=  w8_L2_N5_37;
                        5: B  <=  w8_L2_N6_37;
                        6: B  <=  w8_L2_N7_37;
                        7: B  <=  w8_L2_N8_37;
                        8: B  <=  w8_L2_N9_37;
                        9: B  <= w8_L2_N10_37;
                        10:B  <= w8_L2_N11_37;
                        11:B  <= w8_L2_N12_37;
                        12:B  <= w8_L2_N13_37;
                        13:B  <= w8_L2_N14_37;
                        14:B  <= w8_L2_N15_37;
                        15:B  <= w8_L2_N16_37;
                        16:B  <= w8_L2_N17_37;
                        17:B  <= w8_L2_N18_37;
                        18:B  <= w8_L2_N19_37;
                        19:B  <= w8_L2_N20_37;
                    endcase
                end

               38: begin
                    A  <= N39_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_38;
                        1: B  <=  w8_L2_N2_38;
                        2: B  <=  w8_L2_N3_38;
                        3: B  <=  w8_L2_N4_38;
                        4: B  <=  w8_L2_N5_38;
                        5: B  <=  w8_L2_N6_38;
                        6: B  <=  w8_L2_N7_38;
                        7: B  <=  w8_L2_N8_38;
                        8: B  <=  w8_L2_N9_38;
                        9: B  <= w8_L2_N10_38;
                        10:B  <= w8_L2_N11_38;
                        11:B  <= w8_L2_N12_38;
                        12:B  <= w8_L2_N13_38;
                        13:B  <= w8_L2_N14_38;
                        14:B  <= w8_L2_N15_38;
                        15:B  <= w8_L2_N16_38;
                        16:B  <= w8_L2_N17_38;
                        17:B  <= w8_L2_N18_38;
                        18:B  <= w8_L2_N19_38;
                        19:B  <= w8_L2_N20_38;
                    endcase
                end

               39: begin
                    A  <= N40_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_39;
                        1: B  <=  w8_L2_N2_39;
                        2: B  <=  w8_L2_N3_39;
                        3: B  <=  w8_L2_N4_39;
                        4: B  <=  w8_L2_N5_39;
                        5: B  <=  w8_L2_N6_39;
                        6: B  <=  w8_L2_N7_39;
                        7: B  <=  w8_L2_N8_39;
                        8: B  <=  w8_L2_N9_39;
                        9: B  <= w8_L2_N10_39;
                        10:B  <= w8_L2_N11_39;
                        11:B  <= w8_L2_N12_39;
                        12:B  <= w8_L2_N13_39;
                        13:B  <= w8_L2_N14_39;
                        14:B  <= w8_L2_N15_39;
                        15:B  <= w8_L2_N16_39;
                        16:B  <= w8_L2_N17_39;
                        17:B  <= w8_L2_N18_39;
                        18:B  <= w8_L2_N19_39;
                        19:B  <= w8_L2_N20_39;
                    endcase
                end

               40: begin
                    A  <= N41_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_40;
                        1: B  <=  w8_L2_N2_40;
                        2: B  <=  w8_L2_N3_40;
                        3: B  <=  w8_L2_N4_40;
                        4: B  <=  w8_L2_N5_40;
                        5: B  <=  w8_L2_N6_40;
                        6: B  <=  w8_L2_N7_40;
                        7: B  <=  w8_L2_N8_40;
                        8: B  <=  w8_L2_N9_40;
                        9: B  <= w8_L2_N10_40;
                        10:B  <= w8_L2_N11_40;
                        11:B  <= w8_L2_N12_40;
                        12:B  <= w8_L2_N13_40;
                        13:B  <= w8_L2_N14_40;
                        14:B  <= w8_L2_N15_40;
                        15:B  <= w8_L2_N16_40;
                        16:B  <= w8_L2_N17_40;
                        17:B  <= w8_L2_N18_40;
                        18:B  <= w8_L2_N19_40;
                        19:B  <= w8_L2_N20_40;
                    endcase
                end


               41: begin
                    A  <= N42_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_41;
                        1: B  <=  w8_L2_N2_41;
                        2: B  <=  w8_L2_N3_41;
                        3: B  <=  w8_L2_N4_41;
                        4: B  <=  w8_L2_N5_41;
                        5: B  <=  w8_L2_N6_41;
                        6: B  <=  w8_L2_N7_41;
                        7: B  <=  w8_L2_N8_41;
                        8: B  <=  w8_L2_N9_41;
                        9: B  <= w8_L2_N10_41;
                        10:B  <= w8_L2_N11_41;
                        11:B  <= w8_L2_N12_41;
                        12:B  <= w8_L2_N13_41;
                        13:B  <= w8_L2_N14_41;
                        14:B  <= w8_L2_N15_41;
                        15:B  <= w8_L2_N16_41;
                        16:B  <= w8_L2_N17_41;
                        17:B  <= w8_L2_N18_41;
                        18:B  <= w8_L2_N19_41;
                        19:B  <= w8_L2_N20_41;
                    endcase
                end

               42: begin
                    A  <= N43_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_42;
                        1: B  <=  w8_L2_N2_42;
                        2: B  <=  w8_L2_N3_42;
                        3: B  <=  w8_L2_N4_42;
                        4: B  <=  w8_L2_N5_42;
                        5: B  <=  w8_L2_N6_42;
                        6: B  <=  w8_L2_N7_42;
                        7: B  <=  w8_L2_N8_42;
                        8: B  <=  w8_L2_N9_42;
                        9: B  <= w8_L2_N10_42;
                        10:B  <= w8_L2_N11_42;
                        11:B  <= w8_L2_N12_42;
                        12:B  <= w8_L2_N13_42;
                        13:B  <= w8_L2_N14_42;
                        14:B  <= w8_L2_N15_42;
                        15:B  <= w8_L2_N16_42;
                        16:B  <= w8_L2_N17_42;
                        17:B  <= w8_L2_N18_42;
                        18:B  <= w8_L2_N19_42;
                        19:B  <= w8_L2_N20_42;
                    endcase
                end

               43: begin
                    A  <= N44_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_43;
                        1: B  <=  w8_L2_N2_43;
                        2: B  <=  w8_L2_N3_43;
                        3: B  <=  w8_L2_N4_43;
                        4: B  <=  w8_L2_N5_43;
                        5: B  <=  w8_L2_N6_43;
                        6: B  <=  w8_L2_N7_43;
                        7: B  <=  w8_L2_N8_43;
                        8: B  <=  w8_L2_N9_43;
                        9: B  <= w8_L2_N10_43;
                        10:B  <= w8_L2_N11_43;
                        11:B  <= w8_L2_N12_43;
                        12:B  <= w8_L2_N13_43;
                        13:B  <= w8_L2_N14_43;
                        14:B  <= w8_L2_N15_43;
                        15:B  <= w8_L2_N16_43;
                        16:B  <= w8_L2_N17_43;
                        17:B  <= w8_L2_N18_43;
                        18:B  <= w8_L2_N19_43;
                        19:B  <= w8_L2_N20_43;
                    endcase
                end

               44: begin
                    A  <= N45_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_44;
                        1: B  <=  w8_L2_N2_44;
                        2: B  <=  w8_L2_N3_44;
                        3: B  <=  w8_L2_N4_44;
                        4: B  <=  w8_L2_N5_44;
                        5: B  <=  w8_L2_N6_44;
                        6: B  <=  w8_L2_N7_44;
                        7: B  <=  w8_L2_N8_44;
                        8: B  <=  w8_L2_N9_44;
                        9: B  <= w8_L2_N10_44;
                        10:B  <= w8_L2_N11_44;
                        11:B  <= w8_L2_N12_44;
                        12:B  <= w8_L2_N13_44;
                        13:B  <= w8_L2_N14_44;
                        14:B  <= w8_L2_N15_44;
                        15:B  <= w8_L2_N16_44;
                        16:B  <= w8_L2_N17_44;
                        17:B  <= w8_L2_N18_44;
                        18:B  <= w8_L2_N19_44;
                        19:B  <= w8_L2_N20_44;
                    endcase
                end

               45: begin
                    A  <= N46_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_45;
                        1: B  <=  w8_L2_N2_45;
                        2: B  <=  w8_L2_N3_45;
                        3: B  <=  w8_L2_N4_45;
                        4: B  <=  w8_L2_N5_45;
                        5: B  <=  w8_L2_N6_45;
                        6: B  <=  w8_L2_N7_45;
                        7: B  <=  w8_L2_N8_45;
                        8: B  <=  w8_L2_N9_45;
                        9: B  <= w8_L2_N10_45;
                        10:B  <= w8_L2_N11_45;
                        11:B  <= w8_L2_N12_45;
                        12:B  <= w8_L2_N13_45;
                        13:B  <= w8_L2_N14_45;
                        14:B  <= w8_L2_N15_45;
                        15:B  <= w8_L2_N16_45;
                        16:B  <= w8_L2_N17_45;
                        17:B  <= w8_L2_N18_45;
                        18:B  <= w8_L2_N19_45;
                        19:B  <= w8_L2_N20_45;
                    endcase
                end

               46: begin
                    A  <= N47_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_46;
                        1: B  <=  w8_L2_N2_46;
                        2: B  <=  w8_L2_N3_46;
                        3: B  <=  w8_L2_N4_46;
                        4: B  <=  w8_L2_N5_46;
                        5: B  <=  w8_L2_N6_46;
                        6: B  <=  w8_L2_N7_46;
                        7: B  <=  w8_L2_N8_46;
                        8: B  <=  w8_L2_N9_46;
                        9: B  <= w8_L2_N10_46;
                        10:B  <= w8_L2_N11_46;
                        11:B  <= w8_L2_N12_46;
                        12:B  <= w8_L2_N13_46;
                        13:B  <= w8_L2_N14_46;
                        14:B  <= w8_L2_N15_46;
                        15:B  <= w8_L2_N16_46;
                        16:B  <= w8_L2_N17_46;
                        17:B  <= w8_L2_N18_46;
                        18:B  <= w8_L2_N19_46;
                        19:B  <= w8_L2_N20_46;
                    endcase
                end

               47: begin
                    A  <= N48_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_47;
                        1: B  <=  w8_L2_N2_47;
                        2: B  <=  w8_L2_N3_47;
                        3: B  <=  w8_L2_N4_47;
                        4: B  <=  w8_L2_N5_47;
                        5: B  <=  w8_L2_N6_47;
                        6: B  <=  w8_L2_N7_47;
                        7: B  <=  w8_L2_N8_47;
                        8: B  <=  w8_L2_N9_47;
                        9: B  <= w8_L2_N10_47;
                        10:B  <= w8_L2_N11_47;
                        11:B  <= w8_L2_N12_47;
                        12:B  <= w8_L2_N13_47;
                        13:B  <= w8_L2_N14_47;
                        14:B  <= w8_L2_N15_47;
                        15:B  <= w8_L2_N16_47;
                        16:B  <= w8_L2_N17_47;
                        17:B  <= w8_L2_N18_47;
                        18:B  <= w8_L2_N19_47;
                        19:B  <= w8_L2_N20_47;
                    endcase
                end

               48: begin
                    A  <= N49_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_48;
                        1: B  <=  w8_L2_N2_48;
                        2: B  <=  w8_L2_N3_48;
                        3: B  <=  w8_L2_N4_48;
                        4: B  <=  w8_L2_N5_48;
                        5: B  <=  w8_L2_N6_48;
                        6: B  <=  w8_L2_N7_48;
                        7: B  <=  w8_L2_N8_48;
                        8: B  <=  w8_L2_N9_48;
                        9: B  <= w8_L2_N10_48;
                        10:B  <= w8_L2_N11_48;
                        11:B  <= w8_L2_N12_48;
                        12:B  <= w8_L2_N13_48;
                        13:B  <= w8_L2_N14_48;
                        14:B  <= w8_L2_N15_48;
                        15:B  <= w8_L2_N16_48;
                        16:B  <= w8_L2_N17_48;
                        17:B  <= w8_L2_N18_48;
                        18:B  <= w8_L2_N19_48;
                        19:B  <= w8_L2_N20_48;
                    endcase
                end

               49: begin
                    A  <= N50_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_49;
                        1: B  <=  w8_L2_N2_49;
                        2: B  <=  w8_L2_N3_49;
                        3: B  <=  w8_L2_N4_49;
                        4: B  <=  w8_L2_N5_49;
                        5: B  <=  w8_L2_N6_49;
                        6: B  <=  w8_L2_N7_49;
                        7: B  <=  w8_L2_N8_49;
                        8: B  <=  w8_L2_N9_49;
                        9: B  <= w8_L2_N10_49;
                        10:B  <= w8_L2_N11_49;
                        11:B  <= w8_L2_N12_49;
                        12:B  <= w8_L2_N13_49;
                        13:B  <= w8_L2_N14_49;
                        14:B  <= w8_L2_N15_49;
                        15:B  <= w8_L2_N16_49;
                        16:B  <= w8_L2_N17_49;
                        17:B  <= w8_L2_N18_49;
                        18:B  <= w8_L2_N19_49;
                        19:B  <= w8_L2_N20_49;
                    endcase
                end

               50: begin
                    A  <= N51_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_50;
                        1: B  <=  w8_L2_N2_50;
                        2: B  <=  w8_L2_N3_50;
                        3: B  <=  w8_L2_N4_50;
                        4: B  <=  w8_L2_N5_50;
                        5: B  <=  w8_L2_N6_50;
                        6: B  <=  w8_L2_N7_50;
                        7: B  <=  w8_L2_N8_50;
                        8: B  <=  w8_L2_N9_50;
                        9: B  <= w8_L2_N10_50;
                        10:B  <= w8_L2_N11_50;
                        11:B  <= w8_L2_N12_50;
                        12:B  <= w8_L2_N13_50;
                        13:B  <= w8_L2_N14_50;
                        14:B  <= w8_L2_N15_50;
                        15:B  <= w8_L2_N16_50;
                        16:B  <= w8_L2_N17_50;
                        17:B  <= w8_L2_N18_50;
                        18:B  <= w8_L2_N19_50;
                        19:B  <= w8_L2_N20_50;
                    endcase
                end


               51: begin
                    A  <= N52_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_51;
                        1: B  <=  w8_L2_N2_51;
                        2: B  <=  w8_L2_N3_51;
                        3: B  <=  w8_L2_N4_51;
                        4: B  <=  w8_L2_N5_51;
                        5: B  <=  w8_L2_N6_51;
                        6: B  <=  w8_L2_N7_51;
                        7: B  <=  w8_L2_N8_51;
                        8: B  <=  w8_L2_N9_51;
                        9: B  <= w8_L2_N10_51;
                        10:B  <= w8_L2_N11_51;
                        11:B  <= w8_L2_N12_51;
                        12:B  <= w8_L2_N13_51;
                        13:B  <= w8_L2_N14_51;
                        14:B  <= w8_L2_N15_51;
                        15:B  <= w8_L2_N16_51;
                        16:B  <= w8_L2_N17_51;
                        17:B  <= w8_L2_N18_51;
                        18:B  <= w8_L2_N19_51;
                        19:B  <= w8_L2_N20_51;
                    endcase
                end

               52: begin
                    A  <= N53_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_52;
                        1: B  <=  w8_L2_N2_52;
                        2: B  <=  w8_L2_N3_52;
                        3: B  <=  w8_L2_N4_52;
                        4: B  <=  w8_L2_N5_52;
                        5: B  <=  w8_L2_N6_52;
                        6: B  <=  w8_L2_N7_52;
                        7: B  <=  w8_L2_N8_52;
                        8: B  <=  w8_L2_N9_52;
                        9: B  <= w8_L2_N10_52;
                        10:B  <= w8_L2_N11_52;
                        11:B  <= w8_L2_N12_52;
                        12:B  <= w8_L2_N13_52;
                        13:B  <= w8_L2_N14_52;
                        14:B  <= w8_L2_N15_52;
                        15:B  <= w8_L2_N16_52;
                        16:B  <= w8_L2_N17_52;
                        17:B  <= w8_L2_N18_52;
                        18:B  <= w8_L2_N19_52;
                        19:B  <= w8_L2_N20_52;
                    endcase
                end

               53: begin
                    A  <= N54_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_53;
                        1: B  <=  w8_L2_N2_53;
                        2: B  <=  w8_L2_N3_53;
                        3: B  <=  w8_L2_N4_53;
                        4: B  <=  w8_L2_N5_53;
                        5: B  <=  w8_L2_N6_53;
                        6: B  <=  w8_L2_N7_53;
                        7: B  <=  w8_L2_N8_53;
                        8: B  <=  w8_L2_N9_53;
                        9: B  <= w8_L2_N10_53;
                        10:B  <= w8_L2_N11_53;
                        11:B  <= w8_L2_N12_53;
                        12:B  <= w8_L2_N13_53;
                        13:B  <= w8_L2_N14_53;
                        14:B  <= w8_L2_N15_53;
                        15:B  <= w8_L2_N16_53;
                        16:B  <= w8_L2_N17_53;
                        17:B  <= w8_L2_N18_53;
                        18:B  <= w8_L2_N19_53;
                        19:B  <= w8_L2_N20_53;
                    endcase
                end

               54: begin
                    A  <= N55_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_54;
                        1: B  <=  w8_L2_N2_54;
                        2: B  <=  w8_L2_N3_54;
                        3: B  <=  w8_L2_N4_54;
                        4: B  <=  w8_L2_N5_54;
                        5: B  <=  w8_L2_N6_54;
                        6: B  <=  w8_L2_N7_54;
                        7: B  <=  w8_L2_N8_54;
                        8: B  <=  w8_L2_N9_54;
                        9: B  <= w8_L2_N10_54;
                        10:B  <= w8_L2_N11_54;
                        11:B  <= w8_L2_N12_54;
                        12:B  <= w8_L2_N13_54;
                        13:B  <= w8_L2_N14_54;
                        14:B  <= w8_L2_N15_54;
                        15:B  <= w8_L2_N16_54;
                        16:B  <= w8_L2_N17_54;
                        17:B  <= w8_L2_N18_54;
                        18:B  <= w8_L2_N19_54;
                        19:B  <= w8_L2_N20_54;
                    endcase
                end

               55: begin
                    A  <= N56_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_55;
                        1: B  <=  w8_L2_N2_55;
                        2: B  <=  w8_L2_N3_55;
                        3: B  <=  w8_L2_N4_55;
                        4: B  <=  w8_L2_N5_55;
                        5: B  <=  w8_L2_N6_55;
                        6: B  <=  w8_L2_N7_55;
                        7: B  <=  w8_L2_N8_55;
                        8: B  <=  w8_L2_N9_55;
                        9: B  <= w8_L2_N10_55;
                        10:B  <= w8_L2_N11_55;
                        11:B  <= w8_L2_N12_55;
                        12:B  <= w8_L2_N13_55;
                        13:B  <= w8_L2_N14_55;
                        14:B  <= w8_L2_N15_55;
                        15:B  <= w8_L2_N16_55;
                        16:B  <= w8_L2_N17_55;
                        17:B  <= w8_L2_N18_55;
                        18:B  <= w8_L2_N19_55;
                        19:B  <= w8_L2_N20_55;
                    endcase
                end

               56: begin
                    A  <= N57_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_56;
                        1: B  <=  w8_L2_N2_56;
                        2: B  <=  w8_L2_N3_56;
                        3: B  <=  w8_L2_N4_56;
                        4: B  <=  w8_L2_N5_56;
                        5: B  <=  w8_L2_N6_56;
                        6: B  <=  w8_L2_N7_56;
                        7: B  <=  w8_L2_N8_56;
                        8: B  <=  w8_L2_N9_56;
                        9: B  <= w8_L2_N10_56;
                        10:B  <= w8_L2_N11_56;
                        11:B  <= w8_L2_N12_56;
                        12:B  <= w8_L2_N13_56;
                        13:B  <= w8_L2_N14_56;
                        14:B  <= w8_L2_N15_56;
                        15:B  <= w8_L2_N16_56;
                        16:B  <= w8_L2_N17_56;
                        17:B  <= w8_L2_N18_56;
                        18:B  <= w8_L2_N19_56;
                        19:B  <= w8_L2_N20_56;
                    endcase
                end

               57: begin
                    A  <= N58_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_57;
                        1: B  <=  w8_L2_N2_57;
                        2: B  <=  w8_L2_N3_57;
                        3: B  <=  w8_L2_N4_57;
                        4: B  <=  w8_L2_N5_57;
                        5: B  <=  w8_L2_N6_57;
                        6: B  <=  w8_L2_N7_57;
                        7: B  <=  w8_L2_N8_57;
                        8: B  <=  w8_L2_N9_57;
                        9: B  <= w8_L2_N10_57;
                        10:B  <= w8_L2_N11_57;
                        11:B  <= w8_L2_N12_57;
                        12:B  <= w8_L2_N13_57;
                        13:B  <= w8_L2_N14_57;
                        14:B  <= w8_L2_N15_57;
                        15:B  <= w8_L2_N16_57;
                        16:B  <= w8_L2_N17_57;
                        17:B  <= w8_L2_N18_57;
                        18:B  <= w8_L2_N19_57;
                        19:B  <= w8_L2_N20_57;
                    endcase
                end

               58: begin
                    A  <= N59_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_58;
                        1: B  <=  w8_L2_N2_58;
                        2: B  <=  w8_L2_N3_58;
                        3: B  <=  w8_L2_N4_58;
                        4: B  <=  w8_L2_N5_58;
                        5: B  <=  w8_L2_N6_58;
                        6: B  <=  w8_L2_N7_58;
                        7: B  <=  w8_L2_N8_58;
                        8: B  <=  w8_L2_N9_58;
                        9: B  <= w8_L2_N10_58;
                        10:B  <= w8_L2_N11_58;
                        11:B  <= w8_L2_N12_58;
                        12:B  <= w8_L2_N13_58;
                        13:B  <= w8_L2_N14_58;
                        14:B  <= w8_L2_N15_58;
                        15:B  <= w8_L2_N16_58;
                        16:B  <= w8_L2_N17_58;
                        17:B  <= w8_L2_N18_58;
                        18:B  <= w8_L2_N19_58;
                        19:B  <= w8_L2_N20_58;
                    endcase
                end

               59: begin
                    A  <= N60_L1;
                    C  <= NN_aggre;
                    case(count_NN)
                        0: B  <=  w8_L2_N1_59;
                        1: B  <=  w8_L2_N2_59;
                        2: B  <=  w8_L2_N3_59;
                        3: B  <=  w8_L2_N4_59;
                        4: B  <=  w8_L2_N5_59;
                        5: B  <=  w8_L2_N6_59;
                        6: B  <=  w8_L2_N7_59;
                        7: B  <=  w8_L2_N8_59;
                        8: B  <=  w8_L2_N9_59;
                        9: B  <= w8_L2_N10_59;
                        10:B  <= w8_L2_N11_59;
                        11:B  <= w8_L2_N12_59;
                        12:B  <= w8_L2_N13_59;
                        13:B  <= w8_L2_N14_59;
                        14:B  <= w8_L2_N15_59;
                        15:B  <= w8_L2_N16_59;
                        16:B  <= w8_L2_N17_59;
                        17:B  <= w8_L2_N18_59;
                        18:B  <= w8_L2_N19_59;
                        19:B  <= w8_L2_N20_59;
                    endcase
                end

            endcase
            CE       <= 1;
            count    <= 0;
            nn_state <= waiting_L2_NN;
        end

        waiting_L2_NN: begin
            CE <= 1;
            if(count == 10) begin  //wait done MAC done
                NN_aggre <= P;
                if(count_input == 59)
                    nn_state    <= comp_L2_NN;
                else begin
                    count_input <= count_input + 1; //compute for next input
                    nn_state    <= start_L2_NN;
                end
            end
            else begin
               count    <= count + 1; //wait for MAC operation
               nn_state <= waiting_L2_NN;
            end
        end
        comp_L2_NN: begin
            nn_state    <= next_L2_NN;
            if(NN_aggre[58] == 1)
                NN_aggre <= 59'd0;
        end
        
        next_L2_NN: begin
            if(count_NN == 19) begin
                nn_state    <= done_L2_NN;
                count_input <= 0;
                NN_aggre    <= 0;
                count       <= 0; 
            end  
            else begin
                nn_state    <= start_L2_NN;
                count_NN    <= count_NN + 1;
                count_input <= 0;
                NN_aggre    <= 0;
                count       <= 0;    
            end
            case(count_NN)
                0:  N1_L2  <= NN_aggre[48:19]; //48 --> 10.38    //25 -->  6.19  
                1:  N2_L2  <= NN_aggre[48:19];
                2:  N3_L2  <= NN_aggre[48:19];
                3:  N4_L2  <= NN_aggre[48:19];
                4:  N5_L2  <= NN_aggre[48:19];
                5:  N6_L2  <= NN_aggre[48:19];
                6:  N7_L2  <= NN_aggre[48:19];
                7:  N8_L2  <= NN_aggre[48:19];
                8:  N9_L2  <= NN_aggre[48:19];
                9:  N10_L2 <= NN_aggre[48:19];
                10: N11_L2 <= NN_aggre[48:19]; //48 --> 10.38    //25 -->  6.19  
                11: N12_L2 <= NN_aggre[48:19];
                12: N13_L2 <= NN_aggre[48:19];
                13: N14_L2 <= NN_aggre[48:19];
                14: N15_L2 <= NN_aggre[48:19];
                15: N16_L2 <= NN_aggre[48:19];
                16: N17_L2 <= NN_aggre[48:19];
                17: N18_L2 <= NN_aggre[48:19];
                18: N19_L2 <= NN_aggre[48:19];
                19: N20_L2 <= NN_aggre[48:19];
            endcase
        end
        done_L2_NN: begin
            nn_state    <= start_out_L_NN;   
            count_NN    <= 0;
       end
        start_out_L_NN: begin
                case(count_input)
                    0: begin
                         A  <= N1_L2;
                         case(count_NN)
                             0: begin B  <= w8_out_L_N1_0;   C  <= b_out_L_N1; end
                             1: begin B  <= w8_out_L_N2_0;   C  <= b_out_L_N2; end
                             2: begin B  <= w8_out_L_N3_0;   C  <= b_out_L_N3; end
                        endcase
                    end
                    1: begin
                         A  <= N2_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_1; 
                             1: B  <= w8_out_L_N2_1; 
                             2: B  <= w8_out_L_N3_1; 
                        endcase
                    end
                    2: begin
                         A  <= N3_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_2;
                             1: B  <= w8_out_L_N2_2;
                             2: B  <= w8_out_L_N3_2;
                        endcase
                    end
                    3: begin
                         A  <= N4_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_3;
                             1: B  <= w8_out_L_N2_3;
                             2: B  <= w8_out_L_N3_3;
                        endcase
                    end
                    4: begin
                         A  <= N5_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_4;
                             1: B  <= w8_out_L_N2_4;
                             2: B  <= w8_out_L_N3_4;
                        endcase
                    end
                    5: begin
                         A  <= N6_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_5;
                             1: B  <= w8_out_L_N2_5;
                             2: B  <= w8_out_L_N3_5;
                        endcase
                    end
                    6: begin
                         A  <= N7_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_6;
                             1: B  <= w8_out_L_N2_6;
                             2: B  <= w8_out_L_N3_6;
                        endcase
                    end
                    7: begin
                         A  <= N8_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_7;
                             1: B  <= w8_out_L_N2_7;
                             2: B  <= w8_out_L_N3_7;
                        endcase
                    end
                    8: begin
                         A  <= N9_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_8;
                             1: B  <= w8_out_L_N2_8;
                             2: B  <= w8_out_L_N3_8;
                        endcase
                    end
                    9: begin
                         A  <= N10_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_9;
                             1: B  <= w8_out_L_N2_9;
                             2: B  <= w8_out_L_N3_9;
                        endcase
                    end
                    10: begin
                         A  <= N11_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_10;
                             1: B  <= w8_out_L_N2_10;
                             2: B  <= w8_out_L_N3_10;
                        endcase
                    end
                    11: begin
                         A  <= N12_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_11;
                             1: B  <= w8_out_L_N2_11;
                             2: B  <= w8_out_L_N3_11;
                        endcase
                    end
                    12: begin
                         A  <= N13_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_12;
                             1: B  <= w8_out_L_N2_12;
                             2: B  <= w8_out_L_N3_12;
                        endcase
                    end
                    13: begin
                         A  <= N14_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_13;
                             1: B  <= w8_out_L_N2_13;
                             2: B  <= w8_out_L_N3_13;
                        endcase
                    end
                    14: begin
                         A  <= N15_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_14;
                             1: B  <= w8_out_L_N2_14;
                             2: B  <= w8_out_L_N3_14;
                        endcase
                    end
                    15: begin
                         A  <= N16_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_15;
                             1: B  <= w8_out_L_N2_15;
                             2: B  <= w8_out_L_N3_15;
                        endcase
                    end
                    16: begin
                         A  <= N17_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_16;
                             1: B  <= w8_out_L_N2_16;
                             2: B  <= w8_out_L_N3_16;
                        endcase
                    end
                    17: begin
                         A  <= N18_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_17;
                             1: B  <= w8_out_L_N2_17;
                             2: B  <= w8_out_L_N3_17;
                        endcase
                    end
                    18: begin
                         A  <= N19_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_18;
                             1: B  <= w8_out_L_N2_18;
                             2: B  <= w8_out_L_N3_18;
                        endcase
                    end
                    19: begin
                         A  <= N20_L2;
                         C  <= NN_aggre;
                         case(count_NN)
                             0: B  <= w8_out_L_N1_19;
                             1: B  <= w8_out_L_N2_19;
                             2: B  <= w8_out_L_N3_19;
                        endcase
                    end

                endcase
                CE       <= 1;
                count    <= 0;
                nn_state <= waiting_out_L_NN;
            end   

        waiting_out_L_NN: begin
            CE <= 1;
            if(count == 10) begin  //wait done MAC done
                NN_aggre <= P;
                if(count_input == 19)
                    nn_state    <= next_out_L_NN;
                else begin
                    count_input <= count_input + 1; //compute for next input
                    nn_state    <= start_out_L_NN;
                end
            end
            else begin
               count    <= count + 1; //wait for MAC operation
               nn_state <= waiting_out_L_NN;
            end
        end
        next_out_L_NN: begin
            if(count_NN == 2) begin
                nn_state    <= done_out_L_NN;
                count_input <= 0;
                NN_aggre    <= 0;
                count       <= 0; 
            end  
            else begin
                nn_state    <= start_out_L_NN;
                count_NN    <= count_NN + 1;
                count_input <= 0;
                NN_aggre    <= 0;
                count       <= 0;    
            end
            case(count_NN)
                0:  N1_out_L  <= NN_aggre[48:19]; 
                1:  N2_out_L  <= NN_aggre[48:19];
                2:  N3_out_L  <= NN_aggre[48:19];
            endcase
        end
        done_out_L_NN:
            nn_state    <= compare_outputs;  
            
        compare_outputs: begin
            NN_done <= 1;
            nn_state    <= idle;
            if(($signed(N1_out_L) > $signed(N2_out_L)) && ($signed(N1_out_L) > $signed(N3_out_L))) begin
                EB_LB_HD <= 0;  //EB 
                EB_count    <= EB_count +1;
            end
            else if(($signed(N2_out_L) > $signed(N1_out_L)) && ($signed(N2_out_L) > $signed(N3_out_L))) begin
                EB_LB_HD <= 1;  //HD
                HD_count    <= HD_count +1;
            end
            else if(($signed(N3_out_L) > $signed(N1_out_L)) && ($signed(N3_out_L) > $signed(N2_out_L))) begin
                EB_LB_HD <= 2;  //LB
                LB_count    <= LB_count +1;
            end
            else begin
                EB_LB_HD <= 2;
                //LB_count    <= LB_count +1;
            end
        end  
        
    endcase
end
 
endmodule

