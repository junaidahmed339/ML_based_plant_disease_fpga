`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/18/2022 01:00:40 PM
// Design Name: 
// Module Name: TB_NN
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/10/2022 01:58:34 PM
// Design Name: 
// Module Name: test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TB_NN( );
reg clk=0,reset=0,start_fix_conv=0;
reg [31:0] LBP_161, LBP_156, LBP_137, LBP_136, LBP_132, LBP_128, LBP_125, LBP_43, LBP_38, LBP_32, LBP_25, LBP_19, LBP_14, LBP_7;
reg [31:0]a_bin198 , a_bin199, b_bin208;
reg [2:0]EB_LB_HD = 0;
reg NN_done = 0;

reg clk,reset,start_fix_conv;
wire NN_done;

always begin
#5 clk = ~clk;
end
logic [31:0]data[430][17];
initial begin
data[0][0]=32'h3c9ca18c;	data[0][1]=32'h3d144fe3;	data[0][2]=32'h3f7fa8d6;	data[0][3]=32'h3acc3fdf;	data[0][4]=32'h3af39f9f;	data[0][5]=32'h3a9ff5d4;	data[0][6]=32'h3ae4dd65;	data[0][7]=32'h3b01329b;	data[0][8]=32'h3aa9cdc4;	data[0][9]=32'h3b13a711;	data[0][10]=32'h3acc3fdf;	data[0][11]=32'h3af39f9f;	data[0][12]=32'h3ac4dec2;	data[0][13]=32'h3b03a7c0;	data[0][14]=32'h3a9ff5d4;	data[0][15]=32'h3b01329b;	data[0][16]=32'h3b13a711;
data[1][0]=32'h399302a7;	data[1][1]=32'h00000000;	data[1][2]=32'h3f5e65bf;	data[1][3]=32'h39e41365;	data[1][4]=32'h3a2dc5cb;	data[1][5]=32'h3a53c895;	data[1][6]=32'h3a07c257;	data[1][7]=32'h3abe1148;	data[1][8]=32'h3a07c257;	data[1][9]=32'h3a9ac513;	data[1][10]=32'h39e41365;	data[1][11]=32'h3a2dc5cb;	data[1][12]=32'h398253d8;	data[1][13]=32'h3ad112ad;	data[1][14]=32'h3a53c895;	data[1][15]=32'h3abe1148;	data[1][16]=32'h3a9ac513;
data[2][0]=32'h00000000;	data[2][1]=32'h00000000;	data[2][2]=32'h3f6f6556;	data[2][3]=32'h3a535bdd;	data[2][4]=32'h3a92eb2a;	data[2][5]=32'h3a4e3481;	data[2][6]=32'h39d883e5;	data[2][7]=32'h3a80e0bb;	data[2][8]=32'h3a2a1e4c;	data[2][9]=32'h3a92eb2a;	data[2][10]=32'h3a535bdd;	data[2][11]=32'h3a92eb2a;	data[2][12]=32'h3a060817;	data[2][13]=32'h3a8373bd;	data[2][14]=32'h3a4e3481;	data[2][15]=32'h3a80e0bb;	data[2][16]=32'h3a92eb2a;
data[3][0]=32'h00000000;	data[3][1]=32'h00000000;	data[3][2]=32'h3f6e24dd;	data[3][3]=32'h3a25c0ef;	data[3][4]=32'h39e70c69;	data[3][5]=32'h3a20bb21;	data[3][6]=32'h39a0bb21;	data[3][7]=32'h3a670c69;	data[3][8]=32'h3a2ac6be;	data[3][9]=32'h39d2f530;	data[3][10]=32'h3a25c0ef;	data[3][11]=32'h39e70c69;	data[3][12]=32'h398ca3e8;	data[3][13]=32'h3a02979f;	data[3][14]=32'h3a20bb21;	data[3][15]=32'h3a670c69;	data[3][16]=32'h39d2f530;
data[4][0]=32'h3c6acc92;	data[4][1]=32'h3d3bf940;	data[4][2]=32'h3f7fb741;	data[4][3]=32'h3a6f9422;	data[4][4]=32'h3a9d5d73;	data[4][5]=32'h3a0cedba;	data[4][6]=32'h39bbe7a2;	data[4][7]=32'h3a9d5d73;	data[4][8]=32'h3a49ff68;	data[4][9]=32'h3a98ac34;	data[4][10]=32'h3a6f9422;	data[4][11]=32'h3a9d5d73;	data[4][12]=32'h3a1652e8;	data[4][13]=32'h3aa91bee;	data[4][14]=32'h3a0cedba;	data[4][15]=32'h3a9d5d73;	data[4][16]=32'h3a98ac34;
data[5][0]=32'h3d4c2d6b;	data[5][1]=32'h3d63c537;	data[5][2]=32'h3f7f342f;	data[5][3]=32'h3a63caeb;	data[5][4]=32'h3b20b872;	data[5][5]=32'h3a88ae90;	data[5][6]=32'h3ac7f349;	data[5][7]=32'h3af2fb35;	data[5][8]=32'h3a72fa89;	data[5][9]=32'h3b2850ed;	data[5][10]=32'h3a63caeb;	data[5][11]=32'h3b20b872;	data[5][12]=32'h3aa70d20;	data[5][13]=32'h3ae651d9;	data[5][14]=32'h3a88ae90;	data[5][15]=32'h3af2fb35;	data[5][16]=32'h3b2850ed;
data[6][0]=32'h395c73df;	data[6][1]=32'h00000000;	data[6][2]=32'h3f731077;	data[6][3]=32'h39b45c3e;	data[6][4]=32'h3a1487e2;	data[6][5]=32'h39fea02f;	data[6][6]=32'h3969670c;	data[6][7]=32'h3a8c9321;	data[6][8]=32'h3a81f73c;	data[6][9]=32'h3aa9c058;	data[6][10]=32'h39b45c3e;	data[6][11]=32'h3a1487e2;	data[6][12]=32'h3a696864;	data[6][13]=32'h3a5ecc7f;	data[6][14]=32'h39fea02f;	data[6][15]=32'h3a8c9321;	data[6][16]=32'h3aa9c058;
data[7][0]=32'h00000000;	data[7][1]=32'h00000000;	data[7][2]=32'h3f52e87d;	data[7][3]=32'h3a4a3c7a;	data[7][4]=32'h3aeb0674;	data[7][5]=32'h3a13939b;	data[7][6]=32'h39032d47;	data[7][7]=32'h3a7b6d74;	data[7][8]=32'h39daa222;	data[7][9]=32'h3a9bc771;	data[7][10]=32'h3a4a3c7a;	data[7][11]=32'h3aeb0674;	data[7][12]=32'h3a3f4e09;	data[7][13]=32'h3a190ad3;	data[7][14]=32'h3a13939b;	data[7][15]=32'h3a7b6d74;	data[7][16]=32'h3a9bc771;
data[8][0]=32'h3b18cf6f;	data[8][1]=32'h00000000;	data[8][2]=32'h3f75c3df;	data[8][3]=32'h3aacce2a;	data[8][4]=32'h3ae01b5e;	data[8][5]=32'h3aa4b480;	data[8][6]=32'h3a173510;	data[8][7]=32'h3b02f43c;	data[8][8]=32'h3a94812c;	data[8][9]=32'h3abfb4b6;	data[8][10]=32'h3aacce2a;	data[8][11]=32'h3ae01b5e;	data[8][12]=32'h3aacce2a;	data[8][13]=32'h3b580362;	data[8][14]=32'h3aa4b480;	data[8][15]=32'h3b02f43c;	data[8][16]=32'h3abfb4b6;
data[9][0]=32'h00000000;	data[9][1]=32'h00000000;	data[9][2]=32'h3f71c23b;	data[9][3]=32'h3a9a6069;	data[9][4]=32'h3af9cf64;	data[9][5]=32'h3aa86a17;	data[9][6]=32'h3a91f637;	data[9][7]=32'h3ac74829;	data[9][8]=32'h3a9a6069;	data[9][9]=32'h3af43343;	data[9][10]=32'h3a9a6069;	data[9][11]=32'h3af9cf64;	data[9][12]=32'h3addbf63;	data[9][13]=32'h3b179258;	data[9][14]=32'h3aa86a17;	data[9][15]=32'h3ac74829;	data[9][16]=32'h3af43343;
data[10][0]=32'h3d41908e;	data[10][1]=32'h3d396e16;	data[10][2]=32'h3f7f88b9;	data[10][3]=32'h3a9cd73c;	data[10][4]=32'h3af51414;	data[10][5]=32'h3ac40eb8;	data[10][6]=32'h3a355a95;	data[10][7]=32'h3af7878b;	data[10][8]=32'h3aba40d9;	data[10][9]=32'h3af7878b;	data[10][10]=32'h3a9cd73c;	data[10][11]=32'h3af51414;	data[10][12]=32'h3a8bb250;	data[10][13]=32'h3b0bb0a3;	data[10][14]=32'h3ac40eb8;	data[10][15]=32'h3af7878b;	data[10][16]=32'h3af7878b;
data[11][0]=32'h3c3291b8;	data[11][1]=32'h3c4cd530;	data[11][2]=32'h3f7fd955;	data[11][3]=32'h3a92c2e6;	data[11][4]=32'h3ac3b0c4;	data[11][5]=32'h39fb99bf;	data[11][6]=32'h3ae6a261;	data[11][7]=32'h3af49b48;	data[11][8]=32'h3a43b019;	data[11][9]=32'h3b0bc672;	data[11][10]=32'h3a92c2e6;	data[11][11]=32'h3ac3b0c4;	data[11][12]=32'h39fb99bf;	data[11][13]=32'h3ae6a261;	data[11][14]=32'h39fb99bf;	data[11][15]=32'h3af49b48;	data[11][16]=32'h3b0bc672;
data[12][0]=32'h3c9bb279;	data[12][1]=32'h3cb7b289;	data[12][2]=32'h3f7faace;	data[12][3]=32'h3a9e3433;	data[12][4]=32'h3b08a124;	data[12][5]=32'h3a9235f8;	data[12][6]=32'h3b02a206;	data[12][7]=32'h3b2dc825;	data[12][8]=32'h3aac951f;	data[12][9]=32'h3afbaf38;	data[12][10]=32'h3a9e3433;	data[12][11]=32'h3b08a124;	data[12][12]=32'h3a817002;	data[12][13]=32'h3b1d012d;	data[12][14]=32'h3a9235f8;	data[12][15]=32'h3b2dc825;	data[12][16]=32'h3afbaf38;
data[13][0]=32'h3a9c2c1b;	data[13][1]=32'h00000000;	data[13][2]=32'h3f6417ec;	data[13][3]=32'h3a13ad1c;	data[13][4]=32'h3a8bc317;	data[13][5]=32'h3a1e38e6;	data[13][6]=32'h39680f73;	data[13][7]=32'h3a38980c;	data[13][8]=32'h3a38980c;	data[13][9]=32'h3ab5f443;	data[13][10]=32'h3a13ad1c;	data[13][11]=32'h3a8bc317;	data[13][12]=32'h3a6d55ae;	data[13][13]=32'h3a237f21;	data[13][14]=32'h3a1e38e6;	data[13][15]=32'h3a38980c;	data[13][16]=32'h3ab5f443;
data[14][0]=32'h3cb97fe9;	data[14][1]=32'h3d022ee4;	data[14][2]=32'h3f7fbdcf;	data[14][3]=32'h3a778b92;	data[14][4]=32'h3aeba428;	data[14][5]=32'h3a95f5a0;	data[14][6]=32'h3a87ac31;	data[14][7]=32'h3a82e9d5;	data[14][8]=32'h3a854cdb;	data[14][9]=32'h3af9ed97;	data[14][10]=32'h3a778b92;	data[14][11]=32'h3aeba428;	data[14][12]=32'h3aa69e65;	data[14][13]=32'h3a9f79ad;	data[14][14]=32'h3a95f5a0;	data[14][15]=32'h3a82e9d5;	data[14][16]=32'h3af9ed97;
data[15][0]=32'h39945639;	data[15][1]=32'h00000000;	data[15][2]=32'h3f5fbfc6;	data[15][3]=32'h3a170367;	data[15][4]=32'h3a970210;	data[15][5]=32'h3a8c3888;	data[15][6]=32'h3a27315d;	data[15][7]=32'h3a6d4e4d;	data[15][8]=32'h3a0c39e0;	data[15][9]=32'h3a7817d4;	data[15][10]=32'h3a170367;	data[15][11]=32'h3a970210;	data[15][12]=32'h39e284c5;	data[15][13]=32'h3957bbe9;	data[15][14]=32'h3a8c3888;	data[15][15]=32'h3a6d4e4d;	data[15][16]=32'h3a7817d4;
data[16][0]=32'h37d79654;	data[16][1]=32'h00000000;	data[16][2]=32'h3f5c1c82;	data[16][3]=32'h39947d25;	data[16][4]=32'h3a19cac2;	data[16][5]=32'h39fe8d64;	data[16][6]=32'h38fe8d64;	data[16][7]=32'h3a6ea48e;	data[16][8]=32'h3a0f2f88;	data[16][9]=32'h3ab1a7ad;	data[16][10]=32'h39947d25;	data[16][11]=32'h3a19cac2;	data[16][12]=32'h3a81ed2b;	data[16][13]=32'h3a4ed2e1;	data[16][14]=32'h39fe8d64;	data[16][15]=32'h3a6ea48e;	data[16][16]=32'h3ab1a7ad;
data[17][0]=32'h3b5461ed;	data[17][1]=32'h00000000;	data[17][2]=32'h3f76108c;	data[17][3]=32'h3a50f92c;	data[17][4]=32'h3a813c00;	data[17][5]=32'h3a7cf80e;	data[17][6]=32'h38aff378;	data[17][7]=32'h3a4b79e6;	data[17][8]=32'h3a19fb13;	data[17][9]=32'h3a1f7b05;	data[17][10]=32'h3a50f92c;	data[17][11]=32'h3a813c00;	data[17][12]=32'h3a6c78e5;	data[17][13]=32'h3a7cf80e;	data[17][14]=32'h3a7cf80e;	data[17][15]=32'h3a4b79e6;	data[17][16]=32'h3a1f7b05;
data[18][0]=32'h00000000;	data[18][1]=32'h00000000;	data[18][2]=32'h3f791149;	data[18][3]=32'h3a8ace25;	data[18][4]=32'h3a08493a;	data[18][5]=32'h3a540048;	data[18][6]=32'h39bfcf8e;	data[18][7]=32'h3a1c79f4;	data[18][8]=32'h3a30aaad;	data[18][9]=32'h3a540048;	data[18][10]=32'h3a8ace25;	data[18][11]=32'h3a08493a;	data[18][12]=32'h3a033d62;	data[18][13]=32'h3aae246b;	data[18][14]=32'h3a540048;	data[18][15]=32'h3a1c79f4;	data[18][16]=32'h3a540048;
data[19][0]=32'h3ca85879;	data[19][1]=32'h3d8d2d45;	data[19][2]=32'h3f7f14ba;	data[19][3]=32'h3adf662d;	data[19][4]=32'h3afddf94;	data[19][5]=32'h3a5f6784;	data[19][6]=32'h3ac88da3;	data[19][7]=32'h3ac37b14;	data[19][8]=32'h3ad54110;	data[19][9]=32'h3b040259;	data[19][10]=32'h3adf662d;	data[19][11]=32'h3afddf94;	data[19][12]=32'h3a4b17ec;	data[19][13]=32'h3b068d4d;	data[19][14]=32'h3a5f6784;	data[19][15]=32'h3ac37b14;	data[19][16]=32'h3b040259;
data[20][0]=32'h00000000;	data[20][1]=32'h00000000;	data[20][2]=32'h3f64e465;	data[20][3]=32'h3a38010e;	data[20][4]=32'h3a524a0f;	data[20][5]=32'h3a22f995;	data[20][6]=32'h38fc59ad;	data[20][7]=32'h3a8b5101;	data[20][8]=32'h39b2beda;	data[20][9]=32'h39d24963;	data[20][10]=32'h3a38010e;	data[20][11]=32'h3a524a0f;	data[20][12]=32'h39dccdcc;	data[20][13]=32'h3a1875d8;	data[20][14]=32'h3a22f995;	data[20][15]=32'h3a8b5101;	data[20][16]=32'h39d24963;
data[21][0]=32'h3bffd02f;	data[21][1]=32'h00000000;	data[21][2]=32'h3f587208;	data[21][3]=32'h3a270512;	data[21][4]=32'h3a8963c1;	data[21][5]=32'h3a1c3ee5;	data[21][6]=32'h39b72e55;	data[21][7]=32'h3aac6980;	data[21][8]=32'h39c1f5d9;	data[21][9]=32'h3ab1cc96;	data[21][10]=32'h3a270512;	data[21][11]=32'h3a8963c1;	data[21][12]=32'h3a16db23;	data[21][13]=32'h3abc92c3;	data[21][14]=32'h3a1c3ee5;	data[21][15]=32'h3aac6980;	data[21][16]=32'h3ab1cc96;
data[22][0]=32'h3c4a3a4b;	data[22][1]=32'h3cc00fbb;	data[22][2]=32'h3f7fc30d;	data[22][3]=32'h3aa4a05e;	data[22][4]=32'h3b210e02;	data[22][5]=32'h3ab2f3de;	data[22][6]=32'h3ac60964;	data[22][7]=32'h3af35fdf;	data[22][8]=32'h3a833ab3;	data[22][9]=32'h3adde44c;	data[22][10]=32'h3aa4a05e;	data[22][11]=32'h3b210e02;	data[22][12]=32'h3a9fdafc;	data[22][13]=32'h3b0df6ce;	data[22][14]=32'h3ab2f3de;	data[22][15]=32'h3af35fdf;	data[22][16]=32'h3adde44c;
data[23][0]=32'h3cf15e7d;	data[23][1]=32'h3d07d5ed;	data[23][2]=32'h3f7fc99b;	data[23][3]=32'h3a6ec773;	data[23][4]=32'h3a78868f;	data[23][5]=32'h3a650858;	data[23][6]=32'h3a69e7e6;	data[23][7]=32'h3a86020d;	data[23][8]=32'h3a8391f0;	data[23][9]=32'h3a997f98;	data[23][10]=32'h3a6ec773;	data[23][11]=32'h3a78868f;	data[23][12]=32'h3a997f98;	data[23][13]=32'h3a78868f;	data[23][14]=32'h3a650858;	data[23][15]=32'h3a86020d;	data[23][16]=32'h3a997f98;
data[24][0]=32'h3b2ff881;	data[24][1]=32'h00000000;	data[24][2]=32'h3f753c36;	data[24][3]=32'h3a35f9a2;	data[24][4]=32'h3ae379b7;	data[24][5]=32'h3aab4594;	data[24][6]=32'h3a40ae5b;	data[24][7]=32'h3a95de23;	data[24][8]=32'h3a3b53ff;	data[24][9]=32'h3ad617cf;	data[24][10]=32'h3a35f9a2;	data[24][11]=32'h3ae379b7;	data[24][12]=32'h3a9de3ab;	data[24][13]=32'h3ad0bb6f;	data[24][14]=32'h3aab4594;	data[24][15]=32'h3a95de23;	data[24][16]=32'h3ad617cf;
data[25][0]=32'h00000000;	data[25][1]=32'h00000000;	data[25][2]=32'h3f5cc101;	data[25][3]=32'h3a597780;	data[25][4]=32'h3989e74a;	data[25][5]=32'h39b456df;	data[25][6]=32'h39e96056;	data[25][7]=32'h3a19d178;	data[25][8]=32'h39d429e3;	data[25][9]=32'h3a8740d2;	data[25][10]=32'h3a597780;	data[25][11]=32'h3989e74a;	data[25][12]=32'h39b456df;	data[25][13]=32'h3a6412ba;	data[25][14]=32'h39b456df;	data[25][15]=32'h3a19d178;	data[25][16]=32'h3a8740d2;
data[26][0]=32'h00000000;	data[26][1]=32'h00000000;	data[26][2]=32'h3f61389b;	data[26][3]=32'h3a329945;	data[26][4]=32'h3a9a3edb;	data[26][5]=32'h3a5de4f8;	data[26][6]=32'h39a25c8c;	data[26][7]=32'h3a53120b;	data[26][8]=32'h39d87bd8;	data[26][9]=32'h3a78f49e;	data[26][10]=32'h3a329945;	data[26][11]=32'h3a9a3edb;	data[26][12]=32'h39a25c8c;	data[26][13]=32'h3a8497aa;	data[26][14]=32'h3a5de4f8;	data[26][15]=32'h3a53120b;	data[26][16]=32'h3a78f49e;
data[27][0]=32'h3aeb0674;	data[27][1]=32'h00000000;	data[27][2]=32'h3f69984a;	data[27][3]=32'h3a7650d5;	data[27][4]=32'h3aa8ad33;	data[27][5]=32'h3a95eeea;	data[27][6]=32'h3a20a3a4;	data[27][7]=32'h3a9b47f0;	data[27][8]=32'h3a0082c7;	data[27][9]=32'h3a8889a7;	data[27][10]=32'h3a7650d5;	data[27][11]=32'h3aa8ad33;	data[27][12]=32'h3abe17fe;	data[27][13]=32'h3ab60f1b;	data[27][14]=32'h3a95eeea;	data[27][15]=32'h3a9b47f0;	data[27][16]=32'h3a8889a7;
data[28][0]=32'h39fd45e6;	data[28][1]=32'h00000000;	data[28][2]=32'h3f5a1ab5;	data[28][3]=32'h39e41a1b;	data[28][4]=32'h3a3fd0e6;	data[28][5]=32'h3a357212;	data[28][6]=32'h3925e52c;	data[28][7]=32'h3a5eeb5d;	data[28][8]=32'h399b8659;	data[28][9]=32'h3a896066;	data[28][10]=32'h39e41a1b;	data[28][11]=32'h3a3fd0e6;	data[28][12]=32'h3a44ffa4;	data[28][13]=32'h3a59bc9f;	data[28][14]=32'h3a357212;	data[28][15]=32'h3a5eeb5d;	data[28][16]=32'h3a896066;
data[29][0]=32'h00000000;	data[29][1]=32'h00000000;	data[29][2]=32'h3f6b2032;	data[29][3]=32'h3a0ddea5;	data[29][4]=32'h3a985f07;	data[29][5]=32'h393d29c2;	data[29][6]=32'h393d29c2;	data[29][7]=32'h3a47aacf;	data[29][8]=32'h39b2a6b1;	data[29][9]=32'h39bd286a;	data[29][10]=32'h3a0ddea5;	data[29][11]=32'h3a985f07;	data[29][12]=32'h3993202e;	data[29][13]=32'h3a0ddea5;	data[29][14]=32'h393d29c2;	data[29][15]=32'h3a47aacf;	data[29][16]=32'h39bd286a;
data[30][0]=32'h3a924d75;	data[30][1]=32'h00000000;	data[30][2]=32'h3f77c5ac;	data[30][3]=32'h3a6674bf;	data[30][4]=32'h3a954725;	data[30][5]=32'h3ae9127e;	data[30][6]=32'h3a3c8e10;	data[30][7]=32'h3ad18167;	data[30][8]=32'h3a92a80e;	data[30][9]=32'h3b04406c;	data[30][10]=32'h3a6674bf;	data[30][11]=32'h3a954725;	data[30][12]=32'h3a56be3d;	data[30][13]=32'h3b0eb96c;	data[30][14]=32'h3ae9127e;	data[30][15]=32'h3ad18167;	data[30][16]=32'h3b04406c;
data[31][0]=32'h3d8f01fc;	data[31][1]=32'h3ddd1a22;	data[31][2]=32'h3f7e00d2;	data[31][3]=32'h3aab9cd1;	data[31][4]=32'h3afc38cb;	data[31][5]=32'h3acad221;	data[31][6]=32'h3a5a6bc7;	data[31][7]=32'h3b0db70d;	data[31][8]=32'h3ac839c0;	data[31][9]=32'h3aef3832;	data[31][10]=32'h3aab9cd1;	data[31][11]=32'h3afc38cb;	data[31][12]=32'h3a94375a;	data[31][13]=32'h3af9a06a;	data[31][14]=32'h3acad221;	data[31][15]=32'h3b0db70d;	data[31][16]=32'h3aef3832;
data[32][0]=32'h3b019dfa;	data[32][1]=32'h00000000;	data[32][2]=32'h3f6be61d;	data[32][3]=32'h3aa0f17d;	data[32][4]=32'h3a90d901;	data[32][5]=32'h3a837062;	data[32][6]=32'h3a10d855;	data[32][7]=32'h3af1688e;	data[32][8]=32'h3a3665ad;	data[32][9]=32'h3a467d7d;	data[32][10]=32'h3aa0f17d;	data[32][11]=32'h3a90d901;	data[32][12]=32'h3a7c22a6;	data[32][13]=32'h3ad693f6;	data[32][14]=32'h3a837062;	data[32][15]=32'h3af1688e;	data[32][16]=32'h3a467d7d;
data[33][0]=32'h3c8db6a2;	data[33][1]=32'h3c98b0d1;	data[33][2]=32'h3f7fcaea;	data[33][3]=32'h3a5863af;	data[33][4]=32'h3abc2abe;	data[33][5]=32'h3a377623;	data[33][6]=32'h3a83b6d9;	data[33][7]=32'h3acca12e;	data[33][8]=32'h3a61cc38;	data[33][9]=32'h3afe047d;	data[33][10]=32'h3a5863af;	data[33][11]=32'h3abc2abe;	data[33][12]=32'h3a6fe8b1;	data[33][13]=32'h3ae1cc38;	data[33][14]=32'h3a377623;	data[33][15]=32'h3acca12e;	data[33][16]=32'h3afe047d;
data[34][0]=32'h3a3c86af;	data[34][1]=32'h00000000;	data[34][2]=32'h3f5c0443;	data[34][3]=32'h3a698ffc;	data[34][4]=32'h3a6edef0;	data[34][5]=32'h39a9dd34;	data[34][6]=32'h397ecb22;	data[34][7]=32'h3a742de5;	data[34][8]=32'h38fecdd1;	data[34][9]=32'h3a4f0536;	data[34][10]=32'h3a698ffc;	data[34][11]=32'h3a6edef0;	data[34][12]=32'h3a49b642;	data[34][13]=32'h3a248e3f;	data[34][14]=32'h39a9dd34;	data[34][15]=32'h3a742de5;	data[34][16]=32'h3a4f0536;
data[35][0]=32'h3c4154ca;	data[35][1]=32'h3c809d49;	data[35][2]=32'h3f7fe5c9;	data[35][3]=32'h3a4ec41e;	data[35][4]=32'h3ad35a86;	data[35][5]=32'h3a6eedb4;	data[35][6]=32'h3a99ee53;	data[35][7]=32'h3ab3339f;	data[35][8]=32'h3a4ec41e;	data[35][9]=32'h3aa7b4e5;	data[35][10]=32'h3a4ec41e;	data[35][11]=32'h3ad35a86;	data[35][12]=32'h3a535bdd;	data[35][13]=32'h3a99ee53;	data[35][14]=32'h3a6eedb4;	data[35][15]=32'h3ab3339f;	data[35][16]=32'h3aa7b4e5;
data[36][0]=32'h37c0f020;	data[36][1]=32'h00000000;	data[36][2]=32'h3f70aefb;	data[36][3]=32'h3a8c8910;	data[36][4]=32'h3b0022d0;	data[36][5]=32'h3aaada34;	data[36][6]=32'h3a61f5d4;	data[36][7]=32'h3ac3a6b3;	data[36][8]=32'h3a8443c7;	data[36][9]=32'h3b02e375;	data[36][10]=32'h3a8c8910;	data[36][11]=32'h3b0022d0;	data[36][12]=32'h3a978efd;	data[36][13]=32'h3acbe8a1;	data[36][14]=32'h3aaada34;	data[36][15]=32'h3ac3a6b3;	data[36][16]=32'h3b02e375;
data[37][0]=32'h3d041249;	data[37][1]=32'h3db5cd0c;	data[37][2]=32'h3f7ed71f;	data[37][3]=32'h3a98de89;	data[37][4]=32'h3ad9a522;	data[37][5]=32'h3a8be800;	data[37][6]=32'h3a5ed289;	data[37][7]=32'h3aba8e06;	data[37][8]=32'h3aad977d;	data[37][9]=32'h3ae69850;	data[37][10]=32'h3a98de89;	data[37][11]=32'h3ad9a522;	data[37][12]=32'h3ae930b1;	data[37][13]=32'h3abd230c;	data[37][14]=32'h3a8be800;	data[37][15]=32'h3aba8e06;	data[37][16]=32'h3ae69850;
data[38][0]=32'h3c496463;	data[38][1]=32'h3c188cbf;	data[38][2]=32'h3f7feda6;	data[38][3]=32'h39d0e058;	data[38][4]=32'h3ab11765;	data[38][5]=32'h39b5a10c;	data[38][6]=32'h3aaa4690;	data[38][7]=32'h3aa1313e;	data[38][8]=32'h3a35a10c;	data[38][9]=32'h3a9392ef;	data[38][10]=32'h39d0e058;	data[38][11]=32'h3ab11765;	data[38][12]=32'h3a08391f;	data[38][13]=32'h3a4c5559;	data[38][14]=32'h39b5a10c;	data[38][15]=32'h3aa1313e;	data[38][16]=32'h3a9392ef;
data[39][0]=32'h3ca01cd6;	data[39][1]=32'h3ca5742e;	data[39][2]=32'h3f7fde94;	data[39][3]=32'h3a17e63b;	data[39][4]=32'h3a87ca64;	data[39][5]=32'h3a17e63b;	data[39][6]=32'h3a6f5bc3;	data[39][7]=32'h3a7d2b0e;	data[39][8]=32'h3a00e2be;	data[39][9]=32'h3a80e2be;	data[39][10]=32'h3a17e63b;	data[39][11]=32'h3a87ca64;	data[39][12]=32'h3a53bd2c;	data[39][13]=32'h3a4f2369;	data[39][14]=32'h3a17e63b;	data[39][15]=32'h3a7d2b0e;	data[39][16]=32'h3a80e2be;
data[40][0]=32'h3d1e364c;	data[40][1]=32'h3d81af7d;	data[40][2]=32'h3f7f27bb;	data[40][3]=32'h3ad8665e;	data[40][4]=32'h3ad5db69;	data[40][5]=32'h3a86f04a;	data[40][6]=32'h3a5af2aa;	data[40][7]=32'h3a9b4b4b;	data[40][8]=32'h3ab9d8d4;	data[40][9]=32'h3afc09d1;	data[40][10]=32'h3ad8665e;	data[40][11]=32'h3ad5db69;	data[40][12]=32'h3a797f88;	data[40][13]=32'h3ab4c2eb;	data[40][14]=32'h3a86f04a;	data[40][15]=32'h3a9b4b4b;	data[40][16]=32'h3afc09d1;
data[41][0]=32'h3c810e88;	data[41][1]=32'h3d109071;	data[41][2]=32'h3f7fa440;	data[41][3]=32'h3a4736b6;	data[41][4]=32'h3ad83764;	data[41][5]=32'h3aa7a0c3;	data[41][6]=32'h3a96a0c1;	data[41][7]=32'h3ab63404;	data[41][8]=32'h3ae6caa5;	data[41][9]=32'h3adaa781;	data[41][10]=32'h3a4736b6;	data[41][11]=32'h3ad83764;	data[41][12]=32'h3ad0edc4;	data[41][13]=32'h3b06d572;	data[41][14]=32'h3aa7a0c3;	data[41][15]=32'h3ab63404;	data[41][16]=32'h3adaa781;
data[42][0]=32'h38e85d4c;	data[42][1]=32'h00000000;	data[42][2]=32'h3f734784;	data[42][3]=32'h3a8ca08d;	data[42][4]=32'h3ab7117a;	data[42][5]=32'h3a0f465a;	data[42][6]=32'h3a04a91d;	data[42][7]=32'h3ab1c5e0;	data[42][8]=32'h3a599100;	data[42][9]=32'h3a7eb5a8;	data[42][10]=32'h3a8ca08d;	data[42][11]=32'h3ab7117a;	data[42][12]=32'h3aaf1cb9;	data[42][13]=32'h3aa9cdc4;	data[42][14]=32'h3a0f465a;	data[42][15]=32'h3ab1c5e0;	data[42][16]=32'h3a7eb5a8;
data[43][0]=32'h3d2f8df8;	data[43][1]=32'h3cd1b717;	data[43][2]=32'h3f7fdc9c;	data[43][3]=32'h39df058a;	data[43][4]=32'h3a55ba87;	data[43][5]=32'h3a229efc;	data[43][6]=32'h3a719b8e;	data[43][7]=32'h3a1953f9;	data[43][8]=32'h3a0218c9;	data[43][9]=32'h3a51155c;	data[43][10]=32'h39df058a;	data[43][11]=32'h3a55ba87;	data[43][12]=32'h39b9d980;	data[43][13]=32'h3a14ae22;	data[43][14]=32'h3a229efc;	data[43][15]=32'h3a1953f9;	data[43][16]=32'h3a51155c;
data[44][0]=32'h3db06ab1;	data[44][1]=32'h00000000;	data[44][2]=32'h3f63f91e;	data[44][3]=32'h3a0db1af;	data[44][4]=32'h3a8585e6;	data[44][5]=32'h39e4e4c7;	data[44][6]=32'h39443046;	data[44][7]=32'h3ab11e1b;	data[44][8]=32'h39fab035;	data[44][9]=32'h3a2e64d8;	data[44][10]=32'h3a0db1af;	data[44][11]=32'h3a8585e6;	data[44][12]=32'h3a237e75;	data[44][13]=32'h3a189812;	data[44][14]=32'h39e4e4c7;	data[44][15]=32'h3ab11e1b;	data[44][16]=32'h3a2e64d8;
data[45][0]=32'h00000000;	data[45][1]=32'h00000000;	data[45][2]=32'h3f5a0c4a;	data[45][3]=32'h3a3244b6;	data[45][4]=32'h390e9de8;	data[45][5]=32'h39ad2d75;	data[45][6]=32'h38a2f2df;	data[45][7]=32'h39cbbd02;	data[45][8]=32'h39ea4c8f;	data[45][9]=32'h3a22fcf0;	data[45][10]=32'h3a3244b6;	data[45][11]=32'h390e9de8;	data[45][12]=32'h3a0e9d3c;	data[45][13]=32'h3a4bbc57;	data[45][14]=32'h39ad2d75;	data[45][15]=32'h39cbbd02;	data[45][16]=32'h3a22fcf0;
data[46][0]=32'h3c8cdea0;	data[46][1]=32'h3caa326e;	data[46][2]=32'h3f7fc45d;	data[46][3]=32'h3a1813de;	data[46][4]=32'h3ac9fb61;	data[46][5]=32'h3a42d959;	data[46][6]=32'h3af4c031;	data[46][7]=32'h3aeffe2a;	data[46][8]=32'h3a8050c8;	data[46][9]=32'h3aa3f53d;	data[46][10]=32'h3a1813de;	data[46][11]=32'h3ac9fb61;	data[46][12]=32'h3a1cd48d;	data[46][13]=32'h3a9a748b;	data[46][14]=32'h3a42d959;	data[46][15]=32'h3aeffe2a;	data[46][16]=32'h3aa3f53d;
data[47][0]=32'h386a762b;	data[47][1]=32'h00000000;	data[47][2]=32'h3f7dd399;	data[47][3]=32'h39f229d4;	data[47][4]=32'h3a3a478f;	data[47][5]=32'h399e5719;	data[47][6]=32'h38ba3a23;	data[47][7]=32'h39d6395d;	data[47][8]=32'h390266a2;	data[47][9]=32'h398bb657;	data[47][10]=32'h39f229d4;	data[47][11]=32'h3a3a478f;	data[47][12]=32'h3982654b;	data[47][13]=32'h3a070dd1;	data[47][14]=32'h399e5719;	data[47][15]=32'h39d6395d;	data[47][16]=32'h398bb657;
data[48][0]=32'h3abf7bab;	data[48][1]=32'h00000000;	data[48][2]=32'h3f631705;	data[48][3]=32'h38d2d3a2;	data[48][4]=32'h3ae2a2f8;	data[48][5]=32'h39c849db;	data[48][6]=32'h39f273a5;	data[48][7]=32'h3a4849db;	data[48][8]=32'h3a2def67;	data[48][9]=32'h3a33344a;	data[48][10]=32'h38d2d3a2;	data[48][11]=32'h3ae2a2f8;	data[48][12]=32'h3a4d8ebf;	data[48][13]=32'h3a8e4e0c;	data[48][14]=32'h39c849db;	data[48][15]=32'h3a4849db;	data[48][16]=32'h3a33344a;
data[49][0]=32'h3a147bce;	data[49][1]=32'h00000000;	data[49][2]=32'h3f549279;	data[49][3]=32'h39ed8f65;	data[49][4]=32'h39e33b4e;	data[49][5]=32'h39f7e37c;	data[49][6]=32'h3877e224;	data[49][7]=32'h3a58e68c;	data[49][8]=32'h39ce9321;	data[49][9]=32'h3a3f1452;	data[49][10]=32'h39ed8f65;	data[49][11]=32'h39e33b4e;	data[49][12]=32'h39e33b4e;	data[49][13]=32'h3a39ea47;	data[49][14]=32'h39f7e37c;	data[49][15]=32'h3a58e68c;	data[49][16]=32'h3a3f1452;
data[50][0]=32'h3ccdab19;	data[50][1]=32'h3ce4ba95;	data[50][2]=32'h3f7fb2ab;	data[50][3]=32'h3aacc774;	data[50][4]=32'h3b019744;	data[50][5]=32'h3a666148;	data[50][6]=32'h3a9e632d;	data[50][7]=32'h3aacc774;	data[50][8]=32'h3a926197;	data[50][9]=32'h3b172f5c;	data[50][10]=32'h3aacc774;	data[50][11]=32'h3b019744;	data[50][12]=32'h3a926197;	data[50][13]=32'h3afe6271;	data[50][14]=32'h3a666148;	data[50][15]=32'h3aacc774;	data[50][16]=32'h3b172f5c;
data[51][0]=32'h3c8c5005;	data[51][1]=32'h3c2d8a11;	data[51][2]=32'h3f7fe282;	data[51][3]=32'h3a29d277;	data[51][4]=32'h3ac0c481;	data[51][5]=32'h3a89b0ee;	data[51][6]=32'h3a99c2b4;	data[51][7]=32'h3a8bfc22;	data[51][8]=32'h3a1c0de8;	data[51][9]=32'h3a9095e5;	data[51][10]=32'h3a29d277;	data[51][11]=32'h3ac0c481;	data[51][12]=32'h3a53217b;	data[51][13]=32'h3a8765ba;	data[51][14]=32'h3a89b0ee;	data[51][15]=32'h3a8bfc22;	data[51][16]=32'h3a9095e5;
data[52][0]=32'h37cbd7da;	data[52][1]=32'h00000000;	data[52][2]=32'h3f65436c;	data[52][3]=32'h3a1f9deb;	data[52][4]=32'h3a9250d0;	data[52][5]=32'h39ff62cc;	data[52][6]=32'h38aa49eb;	data[52][7]=32'h39ea1ae6;	data[52][8]=32'h3a6f6c8a;	data[52][9]=32'h3aa79a0d;	data[52][10]=32'h3a1f9deb;	data[52][11]=32'h3a9250d0;	data[52][12]=32'h3a1f9deb;	data[52][13]=32'h3a5f76f3;	data[52][14]=32'h39ff62cc;	data[52][15]=32'h39ea1ae6;	data[52][16]=32'h3aa79a0d;
data[53][0]=32'h3a069256;	data[53][1]=32'h00000000;	data[53][2]=32'h3f55dc1e;	data[53][3]=32'h3a9e9c38;	data[53][4]=32'h3a6f3786;	data[53][5]=32'h39c59d59;	data[53][6]=32'h38d00998;	data[53][7]=32'h3aa90471;	data[53][8]=32'h3a4069e8;	data[53][9]=32'h3a6f3786;	data[53][10]=32'h3a9e9c38;	data[53][11]=32'h3a6f3786;	data[53][12]=32'h39873569;	data[53][13]=32'h3a746af6;	data[53][14]=32'h39c59d59;	data[53][15]=32'h3aa90471;	data[53][16]=32'h3a6f3786;
data[54][0]=32'h3cc7e069;	data[54][1]=32'h00000000;	data[54][2]=32'h3f687358;	data[54][3]=32'h39bbe64b;	data[54][4]=32'h3a827c1c;	data[54][5]=32'h3a027c1c;	data[54][6]=32'h39a705be;	data[54][7]=32'h3a2c3d35;	data[54][8]=32'h3a07b43f;	data[54][9]=32'h3a1c94cc;	data[54][10]=32'h39bbe64b;	data[54][11]=32'h3a827c1c;	data[54][12]=32'h39bbe64b;	data[54][13]=32'h3a270512;	data[54][14]=32'h3a027c1c;	data[54][15]=32'h3a2c3d35;	data[54][16]=32'h3a1c94cc;
data[55][0]=32'h3cb7c99b;	data[55][1]=32'h3d17edc8;	data[55][2]=32'h3f7f88b9;	data[55][3]=32'h3aa59c06;	data[55][4]=32'h3b1e30d8;	data[55][5]=32'h3abbda36;	data[55][6]=32'h3ac0cb37;	data[55][7]=32'h3b26d770;	data[55][8]=32'h3b0ba692;	data[55][9]=32'h3b35ac1f;	data[55][10]=32'h3aa59c06;	data[55][11]=32'h3b1e30d8;	data[55][12]=32'h3aaf7e07;	data[55][13]=32'h3b16c757;	data[55][14]=32'h3abbda36;	data[55][15]=32'h3b26d770;	data[55][16]=32'h3b35ac1f;
data[56][0]=32'h37bcbe62;	data[56][1]=32'h00000000;	data[56][2]=32'h3f75273d;	data[56][3]=32'h3a156603;	data[56][4]=32'h3ad5caa2;	data[56][5]=32'h3a344ed2;	data[56][6]=32'h3962abb1;	data[56][7]=32'h3adaf153;	data[56][8]=32'h3a2a0171;	data[56][9]=32'h3ab6e280;	data[56][10]=32'h3a156603;	data[56][11]=32'h3ad5caa2;	data[56][12]=32'h3a5337a0;	data[56][13]=32'h3a72206e;	data[56][14]=32'h3a344ed2;	data[56][15]=32'h3adaf153;	data[56][16]=32'h3ab6e280;
data[57][0]=32'h3a02c949;	data[57][1]=32'h00000000;	data[57][2]=32'h3f7a60d4;	data[57][3]=32'h3a874e3d;	data[57][4]=32'h3acea5eb;	data[57][5]=32'h39a74a31;	data[57][6]=32'h39b12176;	data[57][7]=32'h3a587ddb;	data[57][8]=32'h3a360d18;	data[57][9]=32'h3a62551f;	data[57][10]=32'h3a874e3d;	data[57][11]=32'h3acea5eb;	data[57][12]=32'h39a74a31;	data[57][13]=32'h3a3fe45c;	data[57][14]=32'h39a74a31;	data[57][15]=32'h3a587ddb;	data[57][16]=32'h3a62551f;
data[58][0]=32'h3995a066;	data[58][1]=32'h00000000;	data[58][2]=32'h3f6cfb55;	data[58][3]=32'h3a841828;	data[58][4]=32'h3a9f0e4e;	data[58][5]=32'h3a52455d;	data[58][6]=32'h3a31ec21;	data[58][7]=32'h3a119239;	data[58][8]=32'h3a8165f1;	data[58][9]=32'h3a8165f1;	data[58][10]=32'h3a841828;	data[58][11]=32'h3a9f0e4e;	data[58][12]=32'h3a2c87b3;	data[58][13]=32'h3aca2db6;	data[58][14]=32'h3a52455d;	data[58][15]=32'h3a119239;	data[58][16]=32'h3a8165f1;
data[59][0]=32'h3c5523b3;	data[59][1]=32'h3cdb8dc5;	data[59][2]=32'h3f7fc1be;	data[59][3]=32'h3a928325;	data[59][4]=32'h3abdc0c0;	data[59][5]=32'h3ac026cc;	data[59][6]=32'h3a88e79b;	data[59][7]=32'h3aa823a0;	data[59][8]=32'h3aaa89ac;	data[59][9]=32'h3ae1c8dd;	data[59][10]=32'h3a928325;	data[59][11]=32'h3abdc0c0;	data[59][12]=32'h3ab8f14e;	data[59][13]=32'h3ada935f;	data[59][14]=32'h3ac026cc;	data[59][15]=32'h3aa823a0;	data[59][16]=32'h3ae1c8dd;
data[60][0]=32'h3c2964e9;	data[60][1]=32'h3ccc9c91;	data[60][2]=32'h3f7fbf1f;	data[60][3]=32'h3a78c6fc;	data[60][4]=32'h3aa0465c;	data[60][5]=32'h3a8391f0;	data[60][6]=32'h3a78c6fc;	data[60][7]=32'h3aa0465c;	data[60][8]=32'h3a944ed7;	data[60][9]=32'h3ab10343;	data[60][10]=32'h3a78c6fc;	data[60][11]=32'h3aa0465c;	data[60][12]=32'h3a78c6fc;	data[60][13]=32'h3abcfac8;	data[60][14]=32'h3a8391f0;	data[60][15]=32'h3aa0465c;	data[60][16]=32'h3ab10343;
data[61][0]=32'h3afec065;	data[61][1]=32'h00000000;	data[61][2]=32'h3f6b65aa;	data[61][3]=32'h3a39c965;	data[61][4]=32'h3abf1702;	data[61][5]=32'h3a1f3e9f;	data[61][6]=32'h39f42d39;	data[61][7]=32'h3aa1e66f;	data[61][8]=32'h398a037a;	data[61][9]=32'h3a698f50;	data[61][10]=32'h3a39c965;	data[61][11]=32'h3abf1702;	data[61][12]=32'h3a8f506a;	data[61][13]=32'h3a91f992;	data[61][14]=32'h3a1f3e9f;	data[61][15]=32'h3aa1e66f;	data[61][16]=32'h3a698f50;
data[62][0]=32'h3d0b3b32;	data[62][1]=32'h3d288df3;	data[62][2]=32'h3f7f8d50;	data[62][3]=32'h3afbd421;	data[62][4]=32'h3b388293;	data[62][5]=32'h3ac9f4ab;	data[62][6]=32'h3abd7da4;	data[62][7]=32'h3b3ffcdb;	data[62][8]=32'h3aea5eae;	data[62][9]=32'h3b5a2b5a;	data[62][10]=32'h3afbd421;	data[62][11]=32'h3b388293;	data[62][12]=32'h3aea5eae;	data[62][13]=32'h3b195754;	data[62][14]=32'h3ac9f4ab;	data[62][15]=32'h3b3ffcdb;	data[62][16]=32'h3b5a2b5a;
data[63][0]=32'h38c699ad;	data[63][1]=32'h00000000;	data[63][2]=32'h3f6fdb4d;	data[63][3]=32'h3a182eb5;	data[63][4]=32'h3a9dd2e4;	data[63][5]=32'h3a61744f;	data[63][6]=32'h3a128bde;	data[63][7]=32'h3b0ce8b1;	data[63][8]=32'h3a508bc9;	data[63][9]=32'h3a39ffc1;	data[63][10]=32'h3a182eb5;	data[63][11]=32'h3a9dd2e4;	data[63][12]=32'h3a725cd4;	data[63][13]=32'h3b0ce8b1;	data[63][14]=32'h3a61744f;	data[63][15]=32'h3b0ce8b1;	data[63][16]=32'h3a39ffc1;
data[64][0]=32'h3b818e0a;	data[64][1]=32'h00000000;	data[64][2]=32'h3f6c154d;	data[64][3]=32'h39ef957a;	data[64][4]=32'h3a45ea85;	data[64][5]=32'h39fa0062;	data[64][6]=32'h397a0062;	data[64][7]=32'h3a5abfaa;	data[64][8]=32'h3a11d555;	data[64][9]=32'h3a45ea85;	data[64][10]=32'h39ef957a;	data[64][11]=32'h3a45ea85;	data[64][12]=32'h3a0234f9;	data[64][13]=32'h3a170ac9;	data[64][14]=32'h39fa0062;	data[64][15]=32'h3a5abfaa;	data[64][16]=32'h3a45ea85;
data[65][0]=32'h37c3745e;	data[65][1]=32'h00000000;	data[65][2]=32'h3f6d8f71;	data[65][3]=32'h3a16767a;	data[65][4]=32'h3a93dcc1;	data[65][5]=32'h3a2b377c;	data[65][6]=32'h394f88bf;	data[65][7]=32'h3a54b8d4;	data[65][8]=32'h3a5f1900;	data[65][9]=32'h3aab3828;	data[65][10]=32'h3a16767a;	data[65][11]=32'h3a93dcc1;	data[65][12]=32'h3a6449c1;	data[65][13]=32'h3abac711;	data[65][14]=32'h3a2b377c;	data[65][15]=32'h3a54b8d4;	data[65][16]=32'h3aab3828;
data[66][0]=32'h3ccdcca7;	data[66][1]=32'h3de085b2;	data[66][2]=32'h3f7e4e27;	data[66][3]=32'h3a536542;	data[66][4]=32'h3a82dd15;	data[66][5]=32'h3a586dc0;	data[66][6]=32'h3a353251;	data[66][7]=32'h3ab531a6;	data[66][8]=32'h3a5d763d;	data[66][9]=32'h3a9982f3;	data[66][10]=32'h3a536542;	data[66][11]=32'h3a82dd15;	data[66][12]=32'h3ab02928;	data[66][13]=32'h3a96feb5;	data[66][14]=32'h3a586dc0;	data[66][15]=32'h3ab531a6;	data[66][16]=32'h3a9982f3;
data[67][0]=32'h3d0388ec;	data[67][1]=32'h3d4abe6a;	data[67][2]=32'h3f7f689d;	data[67][3]=32'h3adbecfb;	data[67][4]=32'h3ab171fd;	data[67][5]=32'h3aaef11a;	data[67][6]=32'h3ab8f14e;	data[67][7]=32'h3b1eb207;	data[67][8]=32'h3aca6d77;	data[67][9]=32'h3b06f3a5;	data[67][10]=32'h3adbecfb;	data[67][11]=32'h3ab171fd;	data[67][12]=32'h3a2ef11a;	data[67][13]=32'h3b10f3d9;	data[67][14]=32'h3aaef11a;	data[67][15]=32'h3b1eb207;	data[67][16]=32'h3b06f3a5;
data[68][0]=32'h3be4da0a;	data[68][1]=32'h00000000;	data[68][2]=32'h3f63c212;	data[68][3]=32'h38f6146f;	data[68][4]=32'h3a6bd3ce;	data[68][5]=32'h3a002ade;	data[68][6]=32'h00000000;	data[68][7]=32'h39cd1094;	data[68][8]=32'h39d751e1;	data[68][9]=32'h3a47f09a;	data[68][10]=32'h38f6146f;	data[68][11]=32'h3a6bd3ce;	data[68][12]=32'h39b88f53;	data[68][13]=32'h3823ff4e;	data[68][14]=32'h3a002ade;	data[68][15]=32'h39cd1094;	data[68][16]=32'h3a47f09a;
data[69][0]=32'h37ba3a23;	data[69][1]=32'h00000000;	data[69][2]=32'h3f766e44;	data[69][3]=32'h3a5c05d0;	data[69][4]=32'h3a7fd6e5;	data[69][5]=32'h3a28dad5;	data[69][6]=32'h3a3d52b1;	data[69][7]=32'h3a827a6e;	data[69][8]=32'h3a9e9f93;	data[69][9]=32'h3a8509c0;	data[69][10]=32'h3a5c05d0;	data[69][11]=32'h3a7fd6e5;	data[69][12]=32'h39adf820;	data[69][13]=32'h3af07dac;	data[69][14]=32'h3a28dad5;	data[69][15]=32'h3a827a6e;	data[69][16]=32'h3a8509c0;
data[70][0]=32'h3c07cad0;	data[70][1]=32'h3cb47a5b;	data[70][2]=32'h3f7fee4e;	data[70][3]=32'h3a3ec929;	data[70][4]=32'h3a30d2f1;	data[70][5]=32'h3a30d2f1;	data[70][6]=32'h399e36e2;	data[70][7]=32'h3a5ab441;	data[70][8]=32'h3a1040aa;	data[70][9]=32'h3a68aa79;	data[70][10]=32'h3a3ec929;	data[70][11]=32'h3a30d2f1;	data[70][12]=32'h3a06f24d;	data[70][13]=32'h3a3ec929;	data[70][14]=32'h3a30d2f1;	data[70][15]=32'h3a5ab441;	data[70][16]=32'h3a68aa79;
data[71][0]=32'h3c4a9692;	data[71][1]=32'h3c0a9d7d;	data[71][2]=32'h3f7fec57;	data[71][3]=32'h3a0cbc11;	data[71][4]=32'h3a709c8b;	data[71][5]=32'h39ec1237;	data[71][6]=32'h3a709c8b;	data[71][7]=32'h3a1ee4b2;	data[71][8]=32'h3a114664;	data[71][9]=32'h3a709c8b;	data[71][10]=32'h3a0cbc11;	data[71][11]=32'h3a709c8b;	data[71][12]=32'h39d9e8ea;	data[71][13]=32'h3a3eac4e;	data[71][14]=32'h39ec1237;	data[71][15]=32'h3a1ee4b2;	data[71][16]=32'h3a709c8b;
data[72][0]=32'h3c8096ff;	data[72][1]=32'h3c32bfdb;	data[72][2]=32'h3f7fe910;	data[72][3]=32'h3a17574a;	data[72][4]=32'h3a409d94;	data[72][5]=32'h39c09e40;	data[72][6]=32'h3a3c07d9;	data[72][7]=32'h3a49c9b8;	data[72][8]=32'h3a578b98;	data[72][9]=32'h3a3c07d9;	data[72][10]=32'h3a17574a;	data[72][11]=32'h3a409d94;	data[72][12]=32'h39e54d77;	data[72][13]=32'h3a17574a;	data[72][14]=32'h39c09e40;	data[72][15]=32'h3a49c9b8;	data[72][16]=32'h3a3c07d9;
data[73][0]=32'h3ca06a6e;	data[73][1]=32'h3d1b499d;	data[73][2]=32'h3f7f8fef;	data[73][3]=32'h3a83c7a0;	data[73][4]=32'h3ade1346;	data[73][5]=32'h3a94dbc5;	data[73][6]=32'h3a174de5;	data[73][7]=32'h3ae566f8;	data[73][8]=32'h3aa5f344;	data[73][9]=32'h3adba329;	data[73][10]=32'h3a83c7a0;	data[73][11]=32'h3ade1346;	data[73][12]=32'h3a88a7da;	data[73][13]=32'h3afdcb72;	data[73][14]=32'h3a94dbc5;	data[73][15]=32'h3ae566f8;	data[73][16]=32'h3adba329;
data[74][0]=32'h3c2fc8b0;	data[74][1]=32'h3c6d8905;	data[74][2]=32'h3f7ff0ed;	data[74][3]=32'h3a1f44a9;	data[74][4]=32'h3aa85cab;	data[74][5]=32'h3a1f44a9;	data[74][6]=32'h39eca07d;	data[74][7]=32'h3a483914;	data[74][8]=32'h3a483914;	data[74][9]=32'h3a6ca07d;	data[74][10]=32'h3a1f44a9;	data[74][11]=32'h3aa85cab;	data[74][12]=32'h3a3f1f0f;	data[74][13]=32'h3a712cd3;	data[74][14]=32'h3a1f44a9;	data[74][15]=32'h3a483914;	data[74][16]=32'h3a6ca07d;
data[75][0]=32'h00000000;	data[75][1]=32'h00000000;	data[75][2]=32'h3f67d8ae;	data[75][3]=32'h39baf4b3;	data[75][4]=32'h3a01d456;	data[75][5]=32'h3a11689e;	data[75][6]=32'h399bcc24;	data[75][7]=32'h3a1bcb78;	data[75][8]=32'h3a169a0b;	data[75][9]=32'h38f9447a;	data[75][10]=32'h39baf4b3;	data[75][11]=32'h3a01d456;	data[75][12]=32'h3a3af407;	data[75][13]=32'h3a4556e2;	data[75][14]=32'h3a11689e;	data[75][15]=32'h3a1bcb78;	data[75][16]=32'h38f9447a;
data[76][0]=32'h3c6019b1;	data[76][1]=32'h3c9f6a94;	data[76][2]=32'h3f7fdfe3;	data[76][3]=32'h3a0fa3a2;	data[76][4]=32'h3a222ce6;	data[76][5]=32'h39cbdfe8;	data[76][6]=32'h3a67ad79;	data[76][7]=32'h3a429b9b;	data[76][8]=32'h39d524e0;	data[76][9]=32'h39e7ad79;	data[76][10]=32'h3a0fa3a2;	data[76][11]=32'h3a222ce6;	data[76][12]=32'h3970f119;	data[76][13]=32'h3a67ad79;	data[76][14]=32'h39cbdfe8;	data[76][15]=32'h3a429b9b;	data[76][16]=32'h39e7ad79;
data[77][0]=32'h3c330f8c;	data[77][1]=32'h3c5f5cf2;	data[77][2]=32'h3f7fd36f;	data[77][3]=32'h3a35e62b;	data[77][4]=32'h3a84eee8;	data[77][5]=32'h3a488e4f;	data[77][6]=32'h3a84eee8;	data[77][7]=32'h3ac88da3;	data[77][8]=32'h3a313c4e;	data[77][9]=32'h3a95406f;	data[77][10]=32'h3a35e62b;	data[77][11]=32'h3a84eee8;	data[77][12]=32'h3a3a90b5;	data[77][13]=32'h3acae2e8;	data[77][14]=32'h3a488e4f;	data[77][15]=32'h3ac88da3;	data[77][16]=32'h3a95406f;
data[78][0]=32'h3a33bc86;	data[78][1]=32'h00000000;	data[78][2]=32'h3f57b15b;	data[78][3]=32'h3a2dda99;	data[78][4]=32'h3a747bbd;	data[78][5]=32'h3a490517;	data[78][6]=32'h39c395ec;	data[78][7]=32'h3a4e7396;	data[78][8]=32'h3a181f46;	data[78][9]=32'h3a0d419d;	data[78][10]=32'h3a2dda99;	data[78][11]=32'h3a747bbd;	data[78][12]=32'h3a3349c4;	data[78][13]=32'h3abb6ed6;	data[78][14]=32'h3a490517;	data[78][15]=32'h3a4e7396;	data[78][16]=32'h3a0d419d;
data[79][0]=32'h3938e7e9;	data[79][1]=32'h00000000;	data[79][2]=32'h3f5ad96a;	data[79][3]=32'h39b159d5;	data[79][4]=32'h3a2643cc;	data[79][5]=32'h3aa907cc;	data[79][6]=32'h39ddaf48;	data[79][7]=32'h3a87c709;	data[79][8]=32'h39bc6f32;	data[79][9]=32'h3a15a3c1;	data[79][10]=32'h39b159d5;	data[79][11]=32'h3a2643cc;	data[79][12]=32'h3a92ddbe;	data[79][13]=32'h3aa643cc;	data[79][14]=32'h3aa907cc;	data[79][15]=32'h3a87c709;	data[79][16]=32'h3a15a3c1;
data[80][0]=32'h3cbae254;	data[80][1]=32'h3d1af295;	data[80][2]=32'h3f7f8f47;	data[80][3]=32'h3ad4f088;	data[80][4]=32'h3b1fb613;	data[80][5]=32'h3ae8c1f6;	data[80][6]=32'h3b0be653;	data[80][7]=32'h3b3af2b0;	data[80][8]=32'h3ac890fe;	data[80][9]=32'h3b2722ef;	data[80][10]=32'h3ad4f088;	data[80][11]=32'h3b1fb613;	data[80][12]=32'h3a9491f3;	data[80][13]=32'h3b4ffdda;	data[80][14]=32'h3ae8c1f6;	data[80][15]=32'h3b3af2b0;	data[80][16]=32'h3b2722ef;
data[81][0]=32'h3b95c5d0;	data[81][1]=32'h00000000;	data[81][2]=32'h3f747b89;	data[81][3]=32'h3ab6a61a;	data[81][4]=32'h3adef0bc;	data[81][5]=32'h3abc05d5;	data[81][6]=32'h3a966b11;	data[81][7]=32'h3b2be6a3;	data[81][8]=32'h3a619e96;	data[81][9]=32'h3b0a53ab;	data[81][10]=32'h3ab6a61a;	data[81][11]=32'h3adef0bc;	data[81][12]=32'h3a619e96;	data[81][13]=32'h3b166963;	data[81][14]=32'h3abc05d5;	data[81][15]=32'h3b2be6a3;	data[81][16]=32'h3b0a53ab;
data[82][0]=32'h3b984fed;	data[82][1]=32'h00000000;	data[82][2]=32'h3f485bc0;	data[82][3]=32'h39d6d108;	data[82][4]=32'h3a78bb93;	data[82][5]=32'h3a1e4901;	data[82][6]=32'h39e21ec4;	data[82][7]=32'h3a18a223;	data[82][8]=32'h3a67c64d;	data[82][9]=32'h3a95cd5c;	data[82][10]=32'h39d6d108;	data[82][11]=32'h3a78bb93;	data[82][12]=32'h39ed6dd7;	data[82][13]=32'h3aa11d1c;	data[82][14]=32'h3a1e4901;	data[82][15]=32'h3a18a223;	data[82][16]=32'h3a95cd5c;
data[83][0]=32'h3b950ef0;	data[83][1]=32'h00000000;	data[83][2]=32'h3f5c1e79;	data[83][3]=32'h3a1632b2;	data[83][4]=32'h3a8849e6;	data[83][5]=32'h3a0b1298;	data[83][6]=32'h3990a2a5;	data[83][7]=32'h3a82ba85;	data[83][8]=32'h3974c4e3;	data[83][9]=32'h39bd2463;	data[83][10]=32'h3a1632b2;	data[83][11]=32'h3a8849e6;	data[83][12]=32'h3a0b1298;	data[83][13]=32'h3a82ba85;	data[83][14]=32'h3a0b1298;	data[83][15]=32'h3a82ba85;	data[83][16]=32'h39bd2463;
data[84][0]=32'h3a261e37;	data[84][1]=32'h00000000;	data[84][2]=32'h3f5c562e;	data[84][3]=32'h3a1cf8ca;	data[84][4]=32'h3a178efd;	data[84][5]=32'h3a7e6724;	data[84][6]=32'h39cdb04d;	data[84][7]=32'h3a6e2a6b;	data[84][8]=32'h396e29bf;	data[84][9]=32'h3a9cf8ca;	data[84][10]=32'h3a1cf8ca;	data[84][11]=32'h3a178efd;	data[84][12]=32'h3a73938b;	data[84][13]=32'h3a6e2a6b;	data[84][14]=32'h3a7e6724;	data[84][15]=32'h3a6e2a6b;	data[84][16]=32'h3a9cf8ca;
data[85][0]=32'h37b7b5e4;	data[85][1]=32'h00000000;	data[85][2]=32'h3f76fd22;	data[85][3]=32'h3a249a54;	data[85][4]=32'h3a34085b;	data[85][5]=32'h3a009841;	data[85][6]=32'h3a97bdf7;	data[85][7]=32'h3a9ce14d;	data[85][8]=32'h3a152ba1;	data[85][9]=32'h3a2ee3ae;	data[85][10]=32'h3a249a54;	data[85][11]=32'h3a34085b;	data[85][12]=32'h39ec9dce;	data[85][13]=32'h3af1c326;	data[85][14]=32'h3a009841;	data[85][15]=32'h3a9ce14d;	data[85][16]=32'h3a2ee3ae;
data[86][0]=32'h3c9e9292;	data[86][1]=32'h3c9988d3;	data[86][2]=32'h3f7fc3b5;	data[86][3]=32'h3a74ce49;	data[86][4]=32'h3a9b5c11;	data[86][5]=32'h3a66ae75;	data[86][6]=32'h3a2010ac;	data[86][7]=32'h3a8ae247;	data[86][8]=32'h3a7e38d6;	data[86][9]=32'h3ab53f12;	data[86][10]=32'h3a74ce49;	data[86][11]=32'h3a9b5c11;	data[86][12]=32'h3a2010ac;	data[86][13]=32'h3a8d3ae7;	data[86][14]=32'h3a66ae75;	data[86][15]=32'h3a8ae247;	data[86][16]=32'h3ab53f12;
data[87][0]=32'h00000000;	data[87][1]=32'h00000000;	data[87][2]=32'h3f6ee243;	data[87][3]=32'h3a4cffce;	data[87][4]=32'h3a14a00b;	data[87][5]=32'h38f5fef5;	data[87][6]=32'h39e18063;	data[87][7]=32'h3a47dfd3;	data[87][8]=32'h39ae409b;	data[87][9]=32'h39f6004d;	data[87][10]=32'h3a4cffce;	data[87][11]=32'h3a14a00b;	data[87][12]=32'h38f5fef5;	data[87][13]=32'h3a002021;	data[87][14]=32'h38f5fef5;	data[87][15]=32'h3a47dfd3;	data[87][16]=32'h39f6004d;
data[88][0]=32'h3c6f62fa;	data[88][1]=32'h3c82d9cf;	data[88][2]=32'h3f7fdf3b;	data[88][3]=32'h3a3d0584;	data[88][4]=32'h3ac1a1f6;	data[88][5]=32'h3a61e710;	data[88][6]=32'h3a8c9d32;	data[88][7]=32'h3a8a4ea3;	data[88][8]=32'h3a4f75f4;	data[88][9]=32'h3aace24c;	data[88][10]=32'h3a3d0584;	data[88][11]=32'h3ac1a1f6;	data[88][12]=32'h3a4f75f4;	data[88][13]=32'h3a463dbc;	data[88][14]=32'h3a61e710;	data[88][15]=32'h3a8a4ea3;	data[88][16]=32'h3aace24c;
data[89][0]=32'h3cdb22d1;	data[89][1]=32'h3d346562;	data[89][2]=32'h3f7f837b;	data[89][3]=32'h3ae368f1;	data[89][4]=32'h3ae0f579;	data[89][5]=32'h3a9a0c86;	data[89][6]=32'h3a2b2b67;	data[89][7]=32'h3b054478;	data[89][8]=32'h3a90455d;	data[89][9]=32'h3aefa391;	data[89][10]=32'h3ae368f1;	data[89][11]=32'h3ae0f579;	data[89][12]=32'h3aab2abc;	data[89][13]=32'h3ab7655c;	data[89][14]=32'h3a9a0c86;	data[89][15]=32'h3b054478;	data[89][16]=32'h3aefa391;
data[90][0]=32'h3c57b203;	data[90][1]=32'h3c5ec5f4;	data[90][2]=32'h3f7fe3d2;	data[90][3]=32'h39c1cd95;	data[90][4]=32'h3a8a6cd6;	data[90][5]=32'h39f92c51;	data[90][6]=32'h3a93aa6c;	data[90][7]=32'h3a66b7da;	data[90][8]=32'h3a05d110;	data[90][9]=32'h3a466ab3;	data[90][10]=32'h39c1cd95;	data[90][11]=32'h3a8a6cd6;	data[90][12]=32'h3a41cd95;	data[90][13]=32'h3a9f3337;	data[90][14]=32'h39f92c51;	data[90][15]=32'h3a66b7da;	data[90][16]=32'h3a466ab3;
data[91][0]=32'h3843745e;	data[91][1]=32'h00000000;	data[91][2]=32'h3f6a2489;	data[91][3]=32'h3a643448;	data[91][4]=32'h3a3c83ff;	data[91][5]=32'h3a417a5e;	data[91][6]=32'h398ae7a5;	data[91][7]=32'h3a2da23a;	data[91][8]=32'h39ee205a;	data[91][9]=32'h398ae7a5;	data[91][10]=32'h3a643448;	data[91][11]=32'h3a3c83ff;	data[91][12]=32'h39e434f3;	data[91][13]=32'h3a378e4c;	data[91][14]=32'h3a417a5e;	data[91][15]=32'h3a2da23a;	data[91][16]=32'h398ae7a5;
data[92][0]=32'h38d31ecb;	data[92][1]=32'h00000000;	data[92][2]=32'h3f68cfc0;	data[92][3]=32'h3a7e5256;	data[92][4]=32'h3ab545c8;	data[92][5]=32'h3a22552a;	data[92][6]=32'h3a329137;	data[92][7]=32'h3a634408;	data[92][8]=32'h3ac01960;	data[92][9]=32'h3aa50863;	data[92][10]=32'h3a7e5256;	data[92][11]=32'h3ab545c8;	data[92][12]=32'h3a634408;	data[92][13]=32'h3aad28c3;	data[92][14]=32'h3a22552a;	data[92][15]=32'h3a634408;	data[92][16]=32'h3aa50863;
data[93][0]=32'h3cb32485;	data[93][1]=32'h3c809f62;	data[93][2]=32'h3f7fe910;	data[93][3]=32'h3a53049f;	data[93][4]=32'h3aa2db62;	data[93][5]=32'h3a12cb9f;	data[93][6]=32'h3ae55ce7;	data[93][7]=32'h3a9e44fa;	data[93][8]=32'h3a454214;	data[93][9]=32'h3aac0831;	data[93][10]=32'h3a53049f;	data[93][11]=32'h3aa2db62;	data[93][12]=32'h3a32e875;	data[93][13]=32'h3aa9bcfd;	data[93][14]=32'h3a12cb9f;	data[93][15]=32'h3a9e44fa;	data[93][16]=32'h3aac0831;
data[94][0]=32'h3cf23cc9;	data[94][1]=32'h3d9ea705;	data[94][2]=32'h3f7eef5f;	data[94][3]=32'h3adb6a1f;	data[94][4]=32'h3b327101;	data[94][5]=32'h3af87c7e;	data[94][6]=32'h3b1e9c38;	data[94][7]=32'h3b5e0e3e;	data[94][8]=32'h3ae8a068;	data[94][9]=32'h3b4e3228;	data[94][10]=32'h3adb6a1f;	data[94][11]=32'h3b327101;	data[94][12]=32'h3ace307a;	data[94][13]=32'h3b3fa74a;	data[94][14]=32'h3af87c7e;	data[94][15]=32'h3b5e0e3e;	data[94][16]=32'h3b4e3228;
data[95][0]=32'h399c2611;	data[95][1]=32'h00000000;	data[95][2]=32'h3f5d6042;	data[95][3]=32'h3a081d9b;	data[95][4]=32'h3a4401f8;	data[95][5]=32'h3a9048b8;	data[95][6]=32'h399873d5;	data[95][7]=32'h3a545786;	data[95][8]=32'h3a081d9b;	data[95][9]=32'h3982ac6d;	data[95][10]=32'h3a081d9b;	data[95][11]=32'h3a4401f8;	data[95][12]=32'h3a13014f;	data[95][13]=32'h3a95b93a;	data[95][14]=32'h3a9048b8;	data[95][15]=32'h3a545786;	data[95][16]=32'h3982ac6d;
data[96][0]=32'h38a50bbe;	data[96][1]=32'h00000000;	data[96][2]=32'h3f5f2086;	data[96][3]=32'h3a239343;	data[96][4]=32'h3aa63660;	data[96][5]=32'h39d31008;	data[96][6]=32'h37a89c6c;	data[96][7]=32'h39fd473e;	data[96][8]=32'h3a62e4bc;	data[96][9]=32'h3a814712;	data[96][10]=32'h3a239343;	data[96][11]=32'h3aa63660;	data[96][12]=32'h3a868efb;	data[96][13]=32'h39fd473e;	data[96][14]=32'h39d31008;	data[96][15]=32'h39fd473e;	data[96][16]=32'h3a814712;
data[97][0]=32'h3cea6c1a;	data[97][1]=32'h3c5edf1e;	data[97][2]=32'h3f7fcaea;	data[97][3]=32'h3a4469fd;	data[97][4]=32'h3ac46951;	data[97][5]=32'h3a77db6e;	data[97][6]=32'h3a809af0;	data[97][7]=32'h3ac2140c;	data[97][8]=32'h3a3fbcc4;	data[97][9]=32'h3ab662fe;	data[97][10]=32'h3a4469fd;	data[97][11]=32'h3ac46951;	data[97][12]=32'h3a65268b;	data[97][13]=32'h3acb6c7a;	data[97][14]=32'h3a77db6e;	data[97][15]=32'h3ac2140c;	data[97][16]=32'h3ab662fe;
data[98][0]=32'h3d1320da;	data[98][1]=32'h3d5c10d8;	data[98][2]=32'h3f7f6b3c;	data[98][3]=32'h3aad14a1;	data[98][4]=32'h3ad22c88;	data[98][5]=32'h3a36f7f9;	data[98][6]=32'h3a0a76e7;	data[98][7]=32'h3ae86ab8;	data[98][8]=32'h3a7c336d;	data[98][9]=32'h3ae5f3e5;	data[98][10]=32'h3aad14a1;	data[98][11]=32'h3ad22c88;	data[98][12]=32'h3a994d43;	data[98][13]=32'h3ad9945b;	data[98][14]=32'h3a36f7f9;	data[98][15]=32'h3ae86ab8;	data[98][16]=32'h3ae5f3e5;
data[99][0]=32'h3a91262e;	data[99][1]=32'h00000000;	data[99][2]=32'h3f6d0481;	data[99][3]=32'h39dd33cd;	data[99][4]=32'h3a28884a;	data[99][5]=32'h3a234412;	data[99][6]=32'h38a89c6c;	data[99][7]=32'h3a28884a;	data[99][8]=32'h3a0e3334;	data[99][9]=32'h3a482243;	data[99][10]=32'h39dd33cd;	data[99][11]=32'h3a28884a;	data[99][12]=32'h39fccd1b;	data[99][13]=32'h3a18bba3;	data[99][14]=32'h3a234412;	data[99][15]=32'h3a28884a;	data[99][16]=32'h3a482243;
data[100][0]=32'h3ce7c287;	data[100][1]=32'h3caf33ca;	data[100][2]=32'h3f7fd955;	data[100][3]=32'h39c3fbee;	data[100][4]=32'h3aa5a617;	data[100][5]=32'h3a3151c7;	data[100][6]=32'h3a6dfac5;	data[100][7]=32'h3a35fc51;	data[100][8]=32'h3a3aa6da;	data[100][9]=32'h3a97a67a;	data[100][10]=32'h39c3fbee;	data[100][11]=32'h3aa5a617;	data[100][12]=32'h3a69503b;	data[100][13]=32'h3a35fc51;	data[100][14]=32'h3a3151c7;	data[100][15]=32'h3a35fc51;	data[100][16]=32'h3a97a67a;
data[101][0]=32'h3c45260f;	data[101][1]=32'h3c780560;	data[101][2]=32'h3f7fef9e;	data[101][3]=32'h3a091ea2;	data[101][4]=32'h3a2daefa;	data[101][5]=32'h39b6d310;	data[101][6]=32'h39e4882a;	data[101][7]=32'h3a248ae4;	data[101][8]=32'h39248ae4;	data[101][9]=32'h3a0db057;	data[101][10]=32'h3a091ea2;	data[101][11]=32'h3a2daefa;	data[101][12]=32'h395b64c0;	data[101][13]=32'h3a36d310;	data[101][14]=32'h39b6d310;	data[101][15]=32'h3a248ae4;	data[101][16]=32'h3a0db057;
data[102][0]=32'h3cae3a3b;	data[102][1]=32'h3d01083e;	data[102][2]=32'h3f7fad6d;	data[102][3]=32'h3ad2a1f9;	data[102][4]=32'h3ade997e;	data[102][5]=32'h3a886ecf;	data[102][6]=32'h3a60fd86;	data[102][7]=32'h3ad03bed;	data[102][8]=32'h3a7db5f9;	data[102][9]=32'h3aea9103;	data[102][10]=32'h3ad2a1f9;	data[102][11]=32'h3ade997e;	data[102][12]=32'h3a7db5f9;	data[102][13]=32'h3ac6aa74;	data[102][14]=32'h3a886ecf;	data[102][15]=32'h3ad03bed;	data[102][16]=32'h3aea9103;
data[103][0]=32'h00000000;	data[103][1]=32'h00000000;	data[103][2]=32'h3f75faec;	data[103][3]=32'h3a6ae841;	data[103][4]=32'h3ad36b4c;	data[103][5]=32'h39fa9156;	data[103][6]=32'h39f02110;	data[103][7]=32'h3a6ae841;	data[103][8]=32'h3aa46e09;	data[103][9]=32'h3abe8a14;	data[103][10]=32'h3a6ae841;	data[103][11]=32'h3ad36b4c;	data[103][12]=32'h3a6ae841;	data[103][13]=32'h3a50cee5;	data[103][14]=32'h39fa9156;	data[103][15]=32'h3a6ae841;	data[103][16]=32'h3abe8a14;
data[104][0]=32'h39990778;	data[104][1]=32'h00000000;	data[104][2]=32'h3f5b3eff;	data[104][3]=32'h3a15cf60;	data[104][4]=32'h3990a554;	data[104][5]=32'h3a10a4a8;	data[104][6]=32'h38f7f79e;	data[104][7]=32'h3a0b79f1;	data[104][8]=32'h3a15cf60;	data[104][9]=32'h39afa2f0;	data[104][10]=32'h3a15cf60;	data[104][11]=32'h3990a554;	data[104][12]=32'h3a2fa39c;	data[104][13]=32'h3a15cf60;	data[104][14]=32'h3a10a4a8;	data[104][15]=32'h3a0b79f1;	data[104][16]=32'h39afa2f0;
data[105][0]=32'h38f4d24f;	data[105][1]=32'h00000000;	data[105][2]=32'h3f4a9e6f;	data[105][3]=32'h3875c945;	data[105][4]=32'h39b86059;	data[105][5]=32'h398f673c;	data[105][6]=32'h00000000;	data[105][7]=32'h39ae21bc;	data[105][8]=32'h39e15977;	data[105][9]=32'h39f5d55a;	data[105][10]=32'h3875c945;	data[105][11]=32'h39b86059;	data[105][12]=32'h38a3c99e;	data[105][13]=32'h3923e476;	data[105][14]=32'h398f673c;	data[105][15]=32'h39ae21bc;	data[105][16]=32'h39f5d55a;
data[106][0]=32'h00000000;	data[106][1]=32'h00000000;	data[106][2]=32'h3f5f1fde;	data[106][3]=32'h39d48680;	data[106][4]=32'h3a6f17fb;	data[106][5]=32'h39f46847;	data[106][6]=32'h3a0a245c;	data[106][7]=32'h3a3f46a7;	data[106][8]=32'h393f4550;	data[106][9]=32'h3a5f27c3;	data[106][10]=32'h39d48680;	data[106][11]=32'h3a6f17fb;	data[106][12]=32'h3a1a1540;	data[106][13]=32'h399f64e0;	data[106][14]=32'h39f46847;	data[106][15]=32'h3a3f46a7;	data[106][16]=32'h3a5f27c3;
data[107][0]=32'h3a9b58b6;	data[107][1]=32'h00000000;	data[107][2]=32'h3f635bd5;	data[107][3]=32'h3986a724;	data[107][4]=32'h3a5984ec;	data[107][5]=32'h39b0165e;	data[107][6]=32'h38cf32d9;	data[107][7]=32'h39c4cd4f;	data[107][8]=32'h394f281c;	data[107][9]=32'h3a3a71d6;	data[107][10]=32'h3986a724;	data[107][11]=32'h3a5984ec;	data[107][12]=32'h39c4cd4f;	data[107][13]=32'h3a690e77;	data[107][14]=32'h39b0165e;	data[107][15]=32'h39c4cd4f;	data[107][16]=32'h3a3a71d6;
data[108][0]=32'h391e688b;	data[108][1]=32'h00000000;	data[108][2]=32'h3f7725c4;	data[108][3]=32'h3a80b26d;	data[108][4]=32'h3abe5e75;	data[108][5]=32'h3a860f79;	data[108][6]=32'h3a0b6bd9;	data[108][7]=32'h3a937817;	data[108][8]=32'h3ab0f5d7;	data[108][9]=32'h3ac3bad5;	data[108][10]=32'h3a80b26d;	data[108][11]=32'h3abe5e75;	data[108][12]=32'h3abbae97;	data[108][13]=32'h3b14ce59;	data[108][14]=32'h3a860f79;	data[108][15]=32'h3a937817;	data[108][16]=32'h3ac3bad5;
data[109][0]=32'h3a54ba2c;	data[109][1]=32'h00000000;	data[109][2]=32'h3f7304ab;	data[109][3]=32'h3abd47f5;	data[109][4]=32'h3a9b1c51;	data[109][5]=32'h3ac2897d;	data[109][6]=32'h3a771d83;	data[109][7]=32'h3aec991b;	data[109][8]=32'h3a32c38c;	data[109][9]=32'h3ab02272;	data[109][10]=32'h3abd47f5;	data[109][11]=32'h3a9b1c51;	data[109][12]=32'h3ac52bef;	data[109][13]=32'h3b037210;	data[109][14]=32'h3ac2897d;	data[109][15]=32'h3aec991b;	data[109][16]=32'h3ab02272;
data[110][0]=32'h39522d34;	data[110][1]=32'h00000000;	data[110][2]=32'h3f75bea1;	data[110][3]=32'h39e0b70f;	data[110][4]=32'h3a51648c;	data[110][5]=32'h3a823baf;	data[110][6]=32'h39c21209;	data[110][7]=32'h3a6aee4b;	data[110][8]=32'h39ada4e9;	data[110][9]=32'h3a4c4944;	data[110][10]=32'h39e0b70f;	data[110][11]=32'h3a51648c;	data[110][12]=32'h39d68080;	data[110][13]=32'h3a823baf;	data[110][14]=32'h3a823baf;	data[110][15]=32'h3a6aee4b;	data[110][16]=32'h3a4c4944;
data[111][0]=32'h3a3a7735;	data[111][1]=32'h00000000;	data[111][2]=32'h3f71057d;	data[111][3]=32'h3a582ca7;	data[111][4]=32'h3b366659;	data[111][5]=32'h3a871be9;	data[111][6]=32'h3981b420;	data[111][7]=32'h3b1e1453;	data[111][8]=32'h3a89cf21;	data[111][9]=32'h3a9cb909;	data[111][10]=32'h3a582ca7;	data[111][11]=32'h3b366659;	data[111][12]=32'h3a81b476;	data[111][13]=32'h3adae08c;	data[111][14]=32'h3a871be9;	data[111][15]=32'h3b1e1453;	data[111][16]=32'h3a9cb909;
data[112][0]=32'h38b9cec3;	data[112][1]=32'h00000000;	data[112][2]=32'h3f755bab;	data[112][3]=32'h3a62cf43;	data[112][4]=32'h3a0d20ba;	data[112][5]=32'h3a173510;	data[112][6]=32'h395dc619;	data[112][7]=32'h3a71eec5;	data[112][8]=32'h3a3572be;	data[112][9]=32'h39bf8714;	data[112][10]=32'h3a62cf43;	data[112][11]=32'h3a0d20ba;	data[112][12]=32'h3a2653e7;	data[112][13]=32'h3a214966;	data[112][14]=32'h3a173510;	data[112][15]=32'h3a71eec5;	data[112][16]=32'h39bf8714;
data[113][0]=32'h39cccac9;	data[113][1]=32'h00000000;	data[113][2]=32'h3f6a2728;	data[113][3]=32'h39d1a19e;	data[113][4]=32'h3a5c1ca1;	data[113][5]=32'h3a084284;	data[113][6]=32'h39dc1ca1;	data[113][7]=32'h3a85a419;	data[113][8]=32'h3a27b43a;	data[113][9]=32'h3a92bc30;	data[113][10]=32'h39d1a19e;	data[113][11]=32'h3a5c1ca1;	data[113][12]=32'h39d1a19e;	data[113][13]=32'h3a12bd87;	data[113][14]=32'h3a084284;	data[113][15]=32'h3a85a419;	data[113][16]=32'h3a92bc30;
data[114][0]=32'h3a2369a7;	data[114][1]=32'h00000000;	data[114][2]=32'h3f755da2;	data[114][3]=32'h3a3ea99e;	data[114][4]=32'h3a89b449;	data[114][5]=32'h3a739f9f;	data[114][6]=32'h39144a24;	data[114][7]=32'h3a78eb39;	data[114][8]=32'h3a81c18c;	data[114][9]=32'h3ab16b47;	data[114][10]=32'h3a3ea99e;	data[114][11]=32'h3a89b449;	data[114][12]=32'h3a8c5a16;	data[114][13]=32'h3aa979e1;	data[114][14]=32'h3a739f9f;	data[114][15]=32'h3a78eb39;	data[114][16]=32'h3ab16b47;
data[115][0]=32'h385bc812;	data[115][1]=32'h00000000;	data[115][2]=32'h3f5e368f;	data[115][3]=32'h3a55817c;	data[115][4]=32'h3a101dc5;	data[115][5]=32'h3a8d73f1;	data[115][6]=32'h3a0ac76f;	data[115][7]=32'h3a602e29;	data[115][8]=32'h3a25771d;	data[115][9]=32'h3ac828f9;	data[115][10]=32'h3a55817c;	data[115][11]=32'h3a101dc5;	data[115][12]=32'h3a8571c4;	data[115][13]=32'h3a602e29;	data[115][14]=32'h3a8d73f1;	data[115][15]=32'h3a602e29;	data[115][16]=32'h3ac828f9;
data[116][0]=32'h3ccd4456;	data[116][1]=32'h3d8d490e;	data[116][2]=32'h3f7f4d16;	data[116][3]=32'h3a323d54;	data[116][4]=32'h3aa36199;	data[116][5]=32'h3a9e7099;	data[116][6]=32'h3aaad023;	data[116][7]=32'h3ab23eac;	data[116][8]=32'h3a4ff21b;	data[116][9]=32'h3aeda58a;	data[116][10]=32'h3a323d54;	data[116][11]=32'h3aa36199;	data[116][12]=32'h3a7c8145;	data[116][13]=32'h3aafc47e;	data[116][14]=32'h3a9e7099;	data[116][15]=32'h3ab23eac;	data[116][16]=32'h3aeda58a;
data[117][0]=32'h3a23852b;	data[117][1]=32'h00000000;	data[117][2]=32'h3f6ab9f5;	data[117][3]=32'h3a349548;	data[117][4]=32'h3a24a668;	data[117][5]=32'h3a59c355;	data[117][6]=32'h3a349548;	data[117][7]=32'h3a646296;	data[117][8]=32'h3ab1ee24;	data[117][9]=32'h3a79a116;	data[117][10]=32'h3a349548;	data[117][11]=32'h3a24a668;	data[117][12]=32'h3a646296;	data[117][13]=32'h3ac1db01;	data[117][14]=32'h3a59c355;	data[117][15]=32'h3a646296;	data[117][16]=32'h3a79a116;
data[118][0]=32'h3cf1c53f;	data[118][1]=32'h3e28240b;	data[118][2]=32'h3f7b630b;	data[118][3]=32'h3aee7239;	data[118][4]=32'h3b1e0a42;	data[118][5]=32'h3ac21767;	data[118][6]=32'h3a0aa1da;	data[118][7]=32'h3aff1448;	data[118][8]=32'h3aa39749;	data[118][9]=32'h3b24f949;	data[118][10]=32'h3aee7239;	data[118][11]=32'h3b1e0a42;	data[118][12]=32'h3acff21b;	data[118][13]=32'h3b15b93a;	data[118][14]=32'h3ac21767;	data[118][15]=32'h3aff1448;	data[118][16]=32'h3b24f949;
data[119][0]=32'h3b73a14d;	data[119][1]=32'h00000000;	data[119][2]=32'h3f6594af;	data[119][3]=32'h3ab20246;	data[119][4]=32'h3ab20246;	data[119][5]=32'h3a67f49b;	data[119][6]=32'h3a0c4096;	data[119][7]=32'h3aed585e;	data[119][8]=32'h3a42323f;	data[119][9]=32'h3a78233d;	data[119][10]=32'h3ab20246;	data[119][11]=32'h3ab20246;	data[119][12]=32'h3ab20246;	data[119][13]=32'h3aba1bf0;	data[119][14]=32'h3a67f49b;	data[119][15]=32'h3aed585e;	data[119][16]=32'h3a78233d;
data[120][0]=32'h3c2e1cde;	data[120][1]=32'h3cb0c671;	data[120][2]=32'h3f7fd2c8;	data[120][3]=32'h3a56db19;	data[120][4]=32'h3a9c7948;	data[120][5]=32'h3a0773d2;	data[120][6]=32'h3aacd185;	data[120][7]=32'h3a7c38cb;	data[120][8]=32'h39f2e1b4;	data[120][9]=32'h3ac8d775;	data[120][10]=32'h3a56db19;	data[120][11]=32'h3a9c7948;	data[120][12]=32'h3a3f805e;	data[120][13]=32'h3a1a22ab;	data[120][14]=32'h3a0773d2;	data[120][15]=32'h3a7c38cb;	data[120][16]=32'h3ac8d775;
data[121][0]=32'h3b985fde;	data[121][1]=32'h00000000;	data[121][2]=32'h3f714467;	data[121][3]=32'h3a97bdf7;	data[121][4]=32'h3ac436fc;	data[121][5]=32'h3a514c63;	data[121][6]=32'h393c5dbf;	data[121][7]=32'h3a5bc360;	data[121][8]=32'h3a2cabf0;	data[121][9]=32'h3ad925a1;	data[121][10]=32'h3a97bdf7;	data[121][11]=32'h3ac436fc;	data[121][12]=32'h3a514c63;	data[121][13]=32'h3ac6d613;	data[121][14]=32'h3a514c63;	data[121][15]=32'h3a5bc360;	data[121][16]=32'h3ad925a1;
data[122][0]=32'h3ca24463;	data[122][1]=32'h3d8bc6a8;	data[122][2]=32'h3f7f2cf9;	data[122][3]=32'h3ab68e9d;	data[122][4]=32'h3b05370c;	data[122][5]=32'h3a5e05da;	data[122][6]=32'h3a406beb;	data[122][7]=32'h3abdf315;	data[122][8]=32'h3a67e480;	data[122][9]=32'h3b05370c;	data[122][10]=32'h3ab68e9d;	data[122][11]=32'h3b05370c;	data[122][12]=32'h3a9b697d;	data[122][13]=32'h3accc2bc;	data[122][14]=32'h3a5e05da;	data[122][15]=32'h3abdf315;	data[122][16]=32'h3b05370c;
data[123][0]=32'h00000000;	data[123][1]=32'h00000000;	data[123][2]=32'h3f54a81a;	data[123][3]=32'h38ad03da;	data[123][4]=32'h39e2fee8;	data[123][5]=32'h3a3d29c2;	data[123][6]=32'h39582f57;	data[123][7]=32'h39f89cb4;	data[123][8]=32'h3917549b;	data[123][9]=32'h3a8c85b5;	data[123][10]=32'h38ad03da;	data[123][11]=32'h39e2fee8;	data[123][12]=32'h3a222381;	data[123][13]=32'h3a1cbbb8;	data[123][14]=32'h3a3d29c2;	data[123][15]=32'h39f89cb4;	data[123][16]=32'h3a8c85b5;
data[124][0]=32'h399b4b4b;	data[124][1]=32'h00000000;	data[124][2]=32'h3f657881;	data[124][3]=32'h3a1c46f3;	data[124][4]=32'h3a74d656;	data[124][5]=32'h3a84d76b;	data[124][6]=32'h3879fb03;	data[124][7]=32'h3a65354e;	data[124][8]=32'h3a023baf;	data[124][9]=32'h3a823b59;	data[124][10]=32'h3a1c46f3;	data[124][11]=32'h3a74d656;	data[124][12]=32'h3a40be77;	data[124][13]=32'h3a9ee2af;	data[124][14]=32'h3a84d76b;	data[124][15]=32'h3a65354e;	data[124][16]=32'h3a823b59;
data[125][0]=32'h3a5a7de5;	data[125][1]=32'h00000000;	data[125][2]=32'h3f6d3847;	data[125][3]=32'h3a47d267;	data[125][4]=32'h3a3d931e;	data[125][5]=32'h39ccf1b6;	data[125][6]=32'h3a3d931e;	data[125][7]=32'h3a669042;	data[125][8]=32'h3a801767;	data[125][9]=32'h3a801767;	data[125][10]=32'h3a47d267;	data[125][11]=32'h3a3d931e;	data[125][12]=32'h3a75ef86;	data[125][13]=32'h3a70cf8b;	data[125][14]=32'h39ccf1b6;	data[125][15]=32'h3a669042;	data[125][16]=32'h3a801767;
data[126][0]=32'h37b60865;	data[126][1]=32'h00000000;	data[126][2]=32'h3f7835bd;	data[126][3]=32'h3a706d91;	data[126][4]=32'h3aa7cc62;	data[126][5]=32'h3a1b4698;	data[126][6]=32'h3a023b03;	data[126][7]=32'h3a84bc93;	data[126][8]=32'h39e668aa;	data[126][9]=32'h3acfddf9;	data[126][10]=32'h3a706d91;	data[126][11]=32'h3aa7cc62;	data[126][12]=32'h3a4358db;	data[126][13]=32'h3ac85b4e;	data[126][14]=32'h3a1b4698;	data[126][15]=32'h3a84bc93;	data[126][16]=32'h3acfddf9;
data[127][0]=32'h3ae7f547;	data[127][1]=32'h00000000;	data[127][2]=32'h3f5b4b73;	data[127][3]=32'h3a199919;	data[127][4]=32'h3a199919;	data[127][5]=32'h39385196;	data[127][6]=32'h00000000;	data[127][7]=32'h3a7ae086;	data[127][8]=32'h3923d70a;	data[127][9]=32'h3a28f501;	data[127][10]=32'h3a199919;	data[127][11]=32'h3a199919;	data[127][12]=32'h3999986d;	data[127][13]=32'h3a0f5bd3;	data[127][14]=32'h39385196;	data[127][15]=32'h3a7ae086;	data[127][16]=32'h3a28f501;
data[128][0]=32'h3bf20a74;	data[128][1]=32'h3c8f9b13;	data[128][2]=32'h3f7fb5f2;	data[128][3]=32'h3a380718;	data[128][4]=32'h3a9246bf;	data[128][5]=32'h39ebedfa;	data[128][6]=32'h3a4ae6ef;	data[128][7]=32'h3a995aaf;	data[128][8]=32'h3a08d780;	data[128][9]=32'h3a841ede;	data[128][10]=32'h3a380718;	data[128][11]=32'h3a9246bf;	data[128][12]=32'h3a206f4c;	data[128][13]=32'h3a96feb5;	data[128][14]=32'h39ebedfa;	data[128][15]=32'h3a995aaf;	data[128][16]=32'h3a841ede;
data[129][0]=32'h3c870111;	data[129][1]=32'h3d026677;	data[129][2]=32'h3f7fc30d;	data[129][3]=32'h3a84eee8;	data[129][4]=32'h3adf2311;	data[129][5]=32'h3aa628f4;	data[129][6]=32'h39e3e1bc;	data[129][7]=32'h3ae8a068;	data[129][8]=32'h3a828e90;	data[129][9]=32'h3ada6465;	data[129][10]=32'h3a84eee8;	data[129][11]=32'h3adf2311;	data[129][12]=32'h3a9f0af3;	data[129][13]=32'h3b0e6c3f;	data[129][14]=32'h3aa628f4;	data[129][15]=32'h3ae8a068;	data[129][16]=32'h3ada6465;
data[130][0]=32'h3ccdca8e;	data[130][1]=32'h3cb3d8e0;	data[130][2]=32'h3f7fcaea;	data[130][3]=32'h3a42e167;	data[130][4]=32'h3ad844d0;	data[130][5]=32'h3a6426dc;	data[130][6]=32'h3a90f734;	data[130][7]=32'h3aeb4990;	data[130][8]=32'h3a8e97de;	data[130][9]=32'h3abbbf5e;	data[130][10]=32'h3a42e167;	data[130][11]=32'h3ad844d0;	data[130][12]=32'h3a1819e8;	data[130][13]=32'h3ac7a2c1;	data[130][14]=32'h3a6426dc;	data[130][15]=32'h3aeb4990;	data[130][16]=32'h3abbbf5e;
data[131][0]=32'h39a0bf28;	data[131][1]=32'h00000000;	data[131][2]=32'h3f5da858;	data[131][3]=32'h3a374a85;	data[131][4]=32'h3aa9691a;	data[131][5]=32'h3a2c2f1d;	data[131][6]=32'h37b1d6a7;	data[131][7]=32'h3a8da2eb;	data[131][8]=32'h3a1b8501;	data[131][9]=32'h3a374a85;	data[131][10]=32'h3a374a85;	data[131][11]=32'h3aa9691a;	data[131][12]=32'h3a47f4a1;	data[131][13]=32'h39c7f3f5;	data[131][14]=32'h3a2c2f1d;	data[131][15]=32'h3a8da2eb;	data[131][16]=32'h3a374a85;
data[132][0]=32'h37c9539c;	data[132][1]=32'h00000000;	data[132][2]=32'h3f65e5f3;	data[132][3]=32'h3aa73c1a;	data[132][4]=32'h3ae9086d;	data[132][5]=32'h3a4adf8d;	data[132][6]=32'h3a0397fb;	data[132][7]=32'h3a9f00e2;	data[132][8]=32'h3ac2a455;	data[132][9]=32'h3aee8300;	data[132][10]=32'h3aa73c1a;	data[132][11]=32'h3ae9086d;	data[132][12]=32'h3a914e71;	data[132][13]=32'h3ab4f1e5;	data[132][14]=32'h3a4adf8d;	data[132][15]=32'h3a9f00e2;	data[132][16]=32'h3aee8300;
data[133][0]=32'h3d137e2c;	data[133][1]=32'h3c6e02a7;	data[133][2]=32'h3f7fbb30;	data[133][3]=32'h3a7edfef;	data[133][4]=32'h3acaf3af;	data[133][5]=32'h3aa9ebf7;	data[133][6]=32'h3a3ccbce;	data[133][7]=32'h3ad91eeb;	data[133][8]=32'h3a5dd589;	data[133][9]=32'h3ac3dfbe;	data[133][10]=32'h3a7edfef;	data[133][11]=32'h3acaf3af;	data[133][12]=32'h3a4183c3;	data[133][13]=32'h3aa078b1;	data[133][14]=32'h3aa9ebf7;	data[133][15]=32'h3ad91eeb;	data[133][16]=32'h3ac3dfbe;
data[134][0]=32'h39e78e9a;	data[134][1]=32'h00000000;	data[134][2]=32'h3f69a9fc;	data[134][3]=32'h3a897b3e;	data[134][4]=32'h3a96f7ff;	data[134][5]=32'h3a21bed7;	data[134][6]=32'h3aa9d47a;	data[134][7]=32'h3a8ee1b0;	data[134][8]=32'h3a729e99;	data[134][9]=32'h3b2317c8;	data[134][10]=32'h3a897b3e;	data[134][11]=32'h3a96f7ff;	data[134][12]=32'h3a841828;	data[134][13]=32'h3b2ddfa2;	data[134][14]=32'h3a21bed7;	data[134][15]=32'h3a8ee1b0;	data[134][16]=32'h3b2317c8;
data[135][0]=32'h3c3927d4;	data[135][1]=32'h3ca30fd0;	data[135][2]=32'h3f7fcaea;	data[135][3]=32'h3abd91c6;	data[135][4]=32'h3b141927;	data[135][5]=32'h3ab1b874;	data[135][6]=32'h3b0f5c29;	data[135][7]=32'h3b270d20;	data[135][8]=32'h3a908bd4;	data[135][9]=32'h3b012381;	data[135][10]=32'h3abd91c6;	data[135][11]=32'h3b141927;	data[135][12]=32'h3ac4ac6d;	data[135][13]=32'h3ac70bc3;	data[135][14]=32'h3ab1b874;	data[135][15]=32'h3b270d20;	data[135][16]=32'h3b012381;
data[136][0]=32'h3c592b80;	data[136][1]=32'h3d153693;	data[136][2]=32'h3f7fb00c;	data[136][3]=32'h3a7384c7;	data[136][4]=32'h3a940505;	data[136][5]=32'h3a834ed4;	data[136][6]=32'h3a91a254;	data[136][7]=32'h3ab30eb6;	data[136][8]=32'h3a521866;	data[136][9]=32'h3a940505;	data[136][10]=32'h3a7384c7;	data[136][11]=32'h3a940505;	data[136][12]=32'h3a43c4e6;	data[136][13]=32'h3a8f3fa4;	data[136][14]=32'h3a834ed4;	data[136][15]=32'h3ab30eb6;	data[136][16]=32'h3a940505;
data[137][0]=32'h3962ec1e;	data[137][1]=32'h00000000;	data[137][2]=32'h3f689a02;	data[137][3]=32'h3a6424d8;	data[137][4]=32'h3a598847;	data[137][5]=32'h3a19dd8c;	data[137][6]=32'h39f40fb2;	data[137][7]=32'h3a6ec169;	data[137][8]=32'h3a29c866;	data[137][9]=32'h3a39b294;	data[137][10]=32'h3a6424d8;	data[137][11]=32'h3a598847;	data[137][12]=32'h3a29c866;	data[137][13]=32'h3ab1bbcf;	data[137][14]=32'h3a19dd8c;	data[137][15]=32'h3a6ec169;	data[137][16]=32'h3a39b294;
data[138][0]=32'h3c87a6bd;	data[138][1]=32'h3c0cf978;	data[138][2]=32'h3f7feef6;	data[138][3]=32'h39fe0b33;	data[138][4]=32'h3a038f41;	data[138][5]=32'h3a3e8811;	data[138][6]=32'h39e2d29e;	data[138][7]=32'h3a2c62ca;	data[138][8]=32'h39ebe5ed;	data[138][9]=32'h3a1a3d83;	data[138][10]=32'h39fe0b33;	data[138][11]=32'h3a038f41;	data[138][12]=32'h39479b60;	data[138][13]=32'h3a4311b8;	data[138][14]=32'h3a3e8811;	data[138][15]=32'h3a2c62ca;	data[138][16]=32'h3a1a3d83;
data[139][0]=32'h3e441355;	data[139][1]=32'h00000000;	data[139][2]=32'h3f6d7f0f;	data[139][3]=32'h3a33410b;	data[139][4]=32'h3a59472f;	data[139][5]=32'h3a92a80e;	data[139][6]=32'h3a0d3ae7;	data[139][7]=32'h3a8d3ae7;	data[139][8]=32'h3a12a965;	data[139][9]=32'h3a7f4d53;	data[139][10]=32'h3a33410b;	data[139][11]=32'h3a59472f;	data[139][12]=32'h3a38af89;	data[139][13]=32'h3a28640d;	data[139][14]=32'h3a92a80e;	data[139][15]=32'h3a8d3ae7;	data[139][16]=32'h3a7f4d53;
data[140][0]=32'h3ddc9c4e;	data[140][1]=32'h00000000;	data[140][2]=32'h3f5bd07d;	data[140][3]=32'h3a38254b;	data[140][4]=32'h3a477dd8;	data[140][5]=32'h3a1456e5;	data[140][6]=32'h39758629;	data[140][7]=32'h39c25fe1;	data[140][8]=32'h39997430;	data[140][9]=32'h3a70698a;	data[140][10]=32'h3a38254b;	data[140][11]=32'h3a477dd8;	data[140][12]=32'h3a0a1c4e;	data[140][13]=32'h39d6d666;	data[140][14]=32'h3a1456e5;	data[140][15]=32'h39c25fe1;	data[140][16]=32'h3a70698a;
data[141][0]=32'h3d482be9;	data[141][1]=32'h00000000;	data[141][2]=32'h3f5835bd;	data[141][3]=32'h39f16487;	data[141][4]=32'h3a182eb5;	data[141][5]=32'h39b26ba3;	data[141][6]=32'h00000000;	data[141][7]=32'h39b26ba3;	data[141][8]=32'h38d1e769;	data[141][9]=32'h3a0dafab;	data[141][10]=32'h39f16487;	data[141][11]=32'h3a182eb5;	data[141][12]=32'h39d1e769;	data[141][13]=32'h39c769b6;	data[141][14]=32'h39b26ba3;	data[141][15]=32'h39b26ba3;	data[141][16]=32'h3a0dafab;
data[142][0]=32'h3adf7398;	data[142][1]=32'h00000000;	data[142][2]=32'h3f6e76c9;	data[142][3]=32'h3ac2c288;	data[142][4]=32'h3a2db301;	data[142][5]=32'h3a1de90a;	data[142][6]=32'h399de90a;	data[142][7]=32'h3ac2c288;	data[142][8]=32'h3a32f68d;	data[142][9]=32'h3ad52cee;	data[142][10]=32'h3ac2c288;	data[142][11]=32'h3a2db301;	data[142][12]=32'h3a80f589;	data[142][13]=32'h3a98a57e;	data[142][14]=32'h3a1de90a;	data[142][15]=32'h3ac2c288;	data[142][16]=32'h3ad52cee;
data[143][0]=32'h3c7e004b;	data[143][1]=32'h3c54e4c9;	data[143][2]=32'h3f7fc84b;	data[143][3]=32'h3aa3146d;	data[143][4]=32'h3a86b73f;	data[143][5]=32'h3a2a2b0c;	data[143][6]=32'h3ad96f72;	data[143][7]=32'h3adbcec8;	data[143][8]=32'h3a9741d1;	data[143][9]=32'h3aa3146d;	data[143][10]=32'h3aa3146d;	data[143][11]=32'h3a86b73f;	data[143][12]=32'h3a9741d1;	data[143][13]=32'h3ae5420f;	data[143][14]=32'h3a2a2b0c;	data[143][15]=32'h3adbcec8;	data[143][16]=32'h3aa3146d;
data[144][0]=32'h3b8e4e0c;	data[144][1]=32'h00000000;	data[144][2]=32'h3f677660;	data[144][3]=32'h39cf8209;	data[144][4]=32'h3a20d1f2;	data[144][5]=32'h39f902b6;	data[144][6]=32'h00000000;	data[144][7]=32'h3a5f12f5;	data[144][8]=32'h39bac1b2;	data[144][9]=32'h393ac30a;	data[144][10]=32'h39cf8209;	data[144][11]=32'h3a20d1f2;	data[144][12]=32'h39e4425f;	data[144][13]=32'h3991425d;	data[144][14]=32'h39f902b6;	data[144][15]=32'h3a5f12f5;	data[144][16]=32'h393ac30a;
data[145][0]=32'h3b5810ce;	data[145][1]=32'h00000000;	data[145][2]=32'h3f5e31f9;	data[145][3]=32'h3a52edce;	data[145][4]=32'h3aa27a13;	data[145][5]=32'h3a9712d7;	data[145][6]=32'h3a7522d7;	data[145][7]=32'h3a94375a;	data[145][8]=32'h3a366d0f;	data[145][9]=32'h3ab94531;	data[145][10]=32'h3a52edce;	data[145][11]=32'h3aa27a13;	data[145][12]=32'h3a7522d7;	data[145][13]=32'h3adb7ae5;	data[145][14]=32'h3a9712d7;	data[145][15]=32'h3a94375a;	data[145][16]=32'h3ab94531;
data[146][0]=32'h3d6a53fc;	data[146][1]=32'h3d4662bb;	data[146][2]=32'h3f7f4b1f;	data[146][3]=32'h3a82c191;	data[146][4]=32'h3ab790fb;	data[146][5]=32'h3a9e69e3;	data[146][6]=32'h3ac19e9b;	data[146][7]=32'h3a8f53c5;	data[146][8]=32'h3a8f53c5;	data[146][9]=32'h3ac927fd;	data[146][10]=32'h3a82c191;	data[146][11]=32'h3ab790fb;	data[146][12]=32'h3a8a4b48;	data[146][13]=32'h3ad84175;	data[146][14]=32'h3a9e69e3;	data[146][15]=32'h3a8f53c5;	data[146][16]=32'h3ac927fd;
data[147][0]=32'h3c910e45;	data[147][1]=32'h3db0025c;	data[147][2]=32'h3f7e9e1b;	data[147][3]=32'h3ab7b5e4;	data[147][4]=32'h3b10e4bf;	data[147][5]=32'h3b0f9a3c;	data[147][6]=32'h39c4a3b3;	data[147][7]=32'h3b21b5c8;	data[147][8]=32'h3b03f4ed;	data[147][9]=32'h3b3b956d;	data[147][10]=32'h3ab7b5e4;	data[147][11]=32'h3b10e4bf;	data[147][12]=32'h3abf7850;	data[147][13]=32'h3adbecfb;	data[147][14]=32'h3b0f9a3c;	data[147][15]=32'h3b21b5c8;	data[147][16]=32'h3b3b956d;
data[148][0]=32'h3c99a416;	data[148][1]=32'h00000000;	data[148][2]=32'h3f5cd0bb;	data[148][3]=32'h3a4ddbeb;	data[148][4]=32'h3a8f1760;	data[148][5]=32'h39a0ab06;	data[148][6]=32'h39aab6a2;	data[148][7]=32'h39e6f6f0;	data[148][8]=32'h3948d571;	data[148][9]=32'h3a39c60a;	data[148][10]=32'h3a4ddbeb;	data[148][11]=32'h3a8f1760;	data[148][12]=32'h39828adf;	data[148][13]=32'h390c9524;	data[148][14]=32'h39a0ab06;	data[148][15]=32'h39e6f6f0;	data[148][16]=32'h3a39c60a;
data[149][0]=32'h3c5e7a74;	data[149][1]=32'h3c05659b;	data[149][2]=32'h3f7ff0ed;	data[149][3]=32'h3a6216b6;	data[149][4]=32'h3a4b7a92;	data[149][5]=32'h3a19bd56;	data[149][6]=32'h39fd387a;	data[149][7]=32'h3a22c897;	data[149][8]=32'h3a34df1a;	data[149][9]=32'h3a5485d4;	data[149][10]=32'h3a6216b6;	data[149][11]=32'h3a4b7a92;	data[149][12]=32'h3a1537b5;	data[149][13]=32'h3a274e38;	data[149][14]=32'h3a19bd56;	data[149][15]=32'h3a22c897;	data[149][16]=32'h3a5485d4;
data[150][0]=32'h3aa1dfb9;	data[150][1]=32'h3f7fff58;	data[150][2]=32'h3b9f1a0c;	data[150][3]=32'h00000000;	data[150][4]=32'h00000000;	data[150][5]=32'h00000000;	data[150][6]=32'h00000000;	data[150][7]=32'h00000000;	data[150][8]=32'h00000000;	data[150][9]=32'h00000000;	data[150][10]=32'h00000000;	data[150][11]=32'h00000000;	data[150][12]=32'h00000000;	data[150][13]=32'h00000000;	data[150][14]=32'h00000000;	data[150][15]=32'h00000000;	data[150][16]=32'h00000000;
data[151][0]=32'h3aceaffc;	data[151][1]=32'h3f7ffeb0;	data[151][2]=32'h3bd3be59;	data[151][3]=32'h00000000;	data[151][4]=32'h00000000;	data[151][5]=32'h00000000;	data[151][6]=32'h00000000;	data[151][7]=32'h00000000;	data[151][8]=32'h00000000;	data[151][9]=32'h00000000;	data[151][10]=32'h00000000;	data[151][11]=32'h00000000;	data[151][12]=32'h00000000;	data[151][13]=32'h00000000;	data[151][14]=32'h00000000;	data[151][15]=32'h00000000;	data[151][16]=32'h00000000;
data[152][0]=32'h3b5013a9;	data[152][1]=32'h3f7ffc11;	data[152][2]=32'h3c24052d;	data[152][3]=32'h00000000;	data[152][4]=32'h00000000;	data[152][5]=32'h00000000;	data[152][6]=32'h00000000;	data[152][7]=32'h00000000;	data[152][8]=32'h00000000;	data[152][9]=32'h00000000;	data[152][10]=32'h00000000;	data[152][11]=32'h00000000;	data[152][12]=32'h00000000;	data[152][13]=32'h00000000;	data[152][14]=32'h00000000;	data[152][15]=32'h00000000;	data[152][16]=32'h00000000;
data[153][0]=32'h3b1fac02;	data[153][1]=32'h3f7ffd61;	data[153][2]=32'h3c0cffc3;	data[153][3]=32'h00000000;	data[153][4]=32'h00000000;	data[153][5]=32'h00000000;	data[153][6]=32'h00000000;	data[153][7]=32'h00000000;	data[153][8]=32'h00000000;	data[153][9]=32'h00000000;	data[153][10]=32'h00000000;	data[153][11]=32'h00000000;	data[153][12]=32'h00000000;	data[153][13]=32'h00000000;	data[153][14]=32'h00000000;	data[153][15]=32'h00000000;	data[153][16]=32'h00000000;
data[154][0]=32'h3b0f73a6;	data[154][1]=32'h3f7ffd61;	data[154][2]=32'h3c02eb01;	data[154][3]=32'h00000000;	data[154][4]=32'h00000000;	data[154][5]=32'h00000000;	data[154][6]=32'h00000000;	data[154][7]=32'h00000000;	data[154][8]=32'h00000000;	data[154][9]=32'h00000000;	data[154][10]=32'h00000000;	data[154][11]=32'h00000000;	data[154][12]=32'h00000000;	data[154][13]=32'h00000000;	data[154][14]=32'h00000000;	data[154][15]=32'h00000000;	data[154][16]=32'h00000000;
data[155][0]=32'h3b4b8900;	data[155][1]=32'h3f7ffb6a;	data[155][2]=32'h3c3c408e;	data[155][3]=32'h00000000;	data[155][4]=32'h00000000;	data[155][5]=32'h00000000;	data[155][6]=32'h00000000;	data[155][7]=32'h00000000;	data[155][8]=32'h00000000;	data[155][9]=32'h00000000;	data[155][10]=32'h00000000;	data[155][11]=32'h00000000;	data[155][12]=32'h00000000;	data[155][13]=32'h00000000;	data[155][14]=32'h00000000;	data[155][15]=32'h00000000;	data[155][16]=32'h00000000;
data[156][0]=32'h399192e5;	data[156][1]=32'h3f08c73b;	data[156][2]=32'h00000000;	data[156][3]=32'h00000000;	data[156][4]=32'h38b0ffe8;	data[156][5]=32'h00000000;	data[156][6]=32'h00000000;	data[156][7]=32'h39137365;	data[156][8]=32'h00000000;	data[156][9]=32'h00000000;	data[156][10]=32'h00000000;	data[156][11]=32'h38b0ffe8;	data[156][12]=32'h37ebb84a;	data[156][13]=32'h00000000;	data[156][14]=32'h00000000;	data[156][15]=32'h39137365;	data[156][16]=32'h00000000;
data[157][0]=32'h3b1cd8e9;	data[157][1]=32'h3f7ffc11;	data[157][2]=32'h3c27fc33;	data[157][3]=32'h00000000;	data[157][4]=32'h00000000;	data[157][5]=32'h00000000;	data[157][6]=32'h00000000;	data[157][7]=32'h00000000;	data[157][8]=32'h00000000;	data[157][9]=32'h00000000;	data[157][10]=32'h00000000;	data[157][11]=32'h00000000;	data[157][12]=32'h00000000;	data[157][13]=32'h00000000;	data[157][14]=32'h00000000;	data[157][15]=32'h00000000;	data[157][16]=32'h00000000;
data[158][0]=32'h3b3fea66;	data[158][1]=32'h3f7ffe09;	data[158][2]=32'h3be925c9;	data[158][3]=32'h00000000;	data[158][4]=32'h37e27e0f;	data[158][5]=32'h00000000;	data[158][6]=32'h00000000;	data[158][7]=32'h37e27e0f;	data[158][8]=32'h38627e0f;	data[158][9]=32'h00000000;	data[158][10]=32'h00000000;	data[158][11]=32'h37e27e0f;	data[158][12]=32'h00000000;	data[158][13]=32'h00000000;	data[158][14]=32'h00000000;	data[158][15]=32'h37e27e0f;	data[158][16]=32'h00000000;
data[159][0]=32'h00000000;	data[159][1]=32'h3f15e3fc;	data[159][2]=32'h00000000;	data[159][3]=32'h39786dba;	data[159][4]=32'h39317355;	data[159][5]=32'h388dfa29;	data[159][6]=32'h380dc479;	data[159][7]=32'h39b17355;	data[159][8]=32'h398df622;	data[159][9]=32'h39786dba;	data[159][10]=32'h39786dba;	data[159][11]=32'h39317355;	data[159][12]=32'h39317355;	data[159][13]=32'h3a0df622;	data[159][14]=32'h388dfa29;	data[159][15]=32'h39b17355;	data[159][16]=32'h39786dba;
data[160][0]=32'h3b096066;	data[160][1]=32'h3f7ffd61;	data[160][2]=32'h3c075056;	data[160][3]=32'h00000000;	data[160][4]=32'h00000000;	data[160][5]=32'h00000000;	data[160][6]=32'h00000000;	data[160][7]=32'h00000000;	data[160][8]=32'h00000000;	data[160][9]=32'h00000000;	data[160][10]=32'h00000000;	data[160][11]=32'h00000000;	data[160][12]=32'h00000000;	data[160][13]=32'h00000000;	data[160][14]=32'h00000000;	data[160][15]=32'h00000000;	data[160][16]=32'h00000000;
data[161][0]=32'h3b23400c;	data[161][1]=32'h3f7ffcb9;	data[161][2]=32'h3c0eb9d7;	data[161][3]=32'h00000000;	data[161][4]=32'h00000000;	data[161][5]=32'h00000000;	data[161][6]=32'h00000000;	data[161][7]=32'h37e27e0f;	data[161][8]=32'h00000000;	data[161][9]=32'h00000000;	data[161][10]=32'h00000000;	data[161][11]=32'h00000000;	data[161][12]=32'h00000000;	data[161][13]=32'h00000000;	data[161][14]=32'h00000000;	data[161][15]=32'h37e27e0f;	data[161][16]=32'h00000000;
data[162][0]=32'h00000000;	data[162][1]=32'h3f148e8a;	data[162][2]=32'h00000000;	data[162][3]=32'h388c825a;	data[162][4]=32'h39d2a4a8;	data[162][5]=32'h380c825a;	data[162][6]=32'h380c825a;	data[162][7]=32'h388c825a;	data[162][8]=32'h39e43244;	data[162][9]=32'h3a03a6be;	data[162][10]=32'h388c825a;	data[162][11]=32'h39d2a4a8;	data[162][12]=32'h39c1170c;	data[162][13]=32'h3975be89;	data[162][14]=32'h380c825a;	data[162][15]=32'h388c825a;	data[162][16]=32'h3a03a6be;
data[163][0]=32'h3b561474;	data[163][1]=32'h3f7ffb6a;	data[163][2]=32'h3c3da943;	data[163][3]=32'h00000000;	data[163][4]=32'h00000000;	data[163][5]=32'h00000000;	data[163][6]=32'h00000000;	data[163][7]=32'h00000000;	data[163][8]=32'h00000000;	data[163][9]=32'h00000000;	data[163][10]=32'h00000000;	data[163][11]=32'h00000000;	data[163][12]=32'h00000000;	data[163][13]=32'h00000000;	data[163][14]=32'h00000000;	data[163][15]=32'h00000000;	data[163][16]=32'h00000000;
data[164][0]=32'h3b1aad96;	data[164][1]=32'h3f7ffcb9;	data[164][2]=32'h3c2a6d26;	data[164][3]=32'h00000000;	data[164][4]=32'h00000000;	data[164][5]=32'h00000000;	data[164][6]=32'h00000000;	data[164][7]=32'h00000000;	data[164][8]=32'h00000000;	data[164][9]=32'h00000000;	data[164][10]=32'h00000000;	data[164][11]=32'h00000000;	data[164][12]=32'h00000000;	data[164][13]=32'h00000000;	data[164][14]=32'h00000000;	data[164][15]=32'h00000000;	data[164][16]=32'h00000000;
data[165][0]=32'h00000000;	data[165][1]=32'h3f057d18;	data[165][2]=32'h00000000;	data[165][3]=32'h00000000;	data[165][4]=32'h00000000;	data[165][5]=32'h38b2e317;	data[165][6]=32'h00000000;	data[165][7]=32'h39d09e93;	data[165][8]=32'h3915035d;	data[165][9]=32'h38ee6cdb;	data[165][10]=32'h00000000;	data[165][11]=32'h00000000;	data[165][12]=32'h00000000;	data[165][13]=32'h39d09e93;	data[165][14]=32'h38b2e317;	data[165][15]=32'h39d09e93;	data[165][16]=32'h38ee6cdb;
data[166][0]=32'h00000000;	data[166][1]=32'h3ee031cf;	data[166][2]=32'h00000000;	data[166][3]=32'h00000000;	data[166][4]=32'h00000000;	data[166][5]=32'h00000000;	data[166][6]=32'h00000000;	data[166][7]=32'h3a154dda;	data[166][8]=32'h00000000;	data[166][9]=32'h38b318c7;	data[166][10]=32'h00000000;	data[166][11]=32'h00000000;	data[166][12]=32'h00000000;	data[166][13]=32'h39154e86;	data[166][14]=32'h00000000;	data[166][15]=32'h3a154dda;	data[166][16]=32'h38b318c7;
data[167][0]=32'h3b392550;	data[167][1]=32'h3f7ffc11;	data[167][2]=32'h3c2f965b;	data[167][3]=32'h37e1a74f;	data[167][4]=32'h00000000;	data[167][5]=32'h00000000;	data[167][6]=32'h37e1a74f;	data[167][7]=32'h00000000;	data[167][8]=32'h00000000;	data[167][9]=32'h00000000;	data[167][10]=32'h37e1a74f;	data[167][11]=32'h00000000;	data[167][12]=32'h00000000;	data[167][13]=32'h00000000;	data[167][14]=32'h00000000;	data[167][15]=32'h00000000;	data[167][16]=32'h00000000;
data[168][0]=32'h3b770b65;	data[168][1]=32'h3f7ff823;	data[168][2]=32'h3c7709b7;	data[168][3]=32'h00000000;	data[168][4]=32'h00000000;	data[168][5]=32'h00000000;	data[168][6]=32'h37e27e0f;	data[168][7]=32'h00000000;	data[168][8]=32'h00000000;	data[168][9]=32'h00000000;	data[168][10]=32'h00000000;	data[168][11]=32'h00000000;	data[168][12]=32'h00000000;	data[168][13]=32'h00000000;	data[168][14]=32'h00000000;	data[168][15]=32'h00000000;	data[168][16]=32'h00000000;
data[169][0]=32'h00000000;	data[169][1]=32'h3ef657fb;	data[169][2]=32'h00000000;	data[169][3]=32'h38b2e317;	data[169][4]=32'h3a0da240;	data[169][5]=32'h00000000;	data[169][6]=32'h00000000;	data[169][7]=32'h37ee3c89;	data[169][8]=32'h00000000;	data[169][9]=32'h38ee87b3;	data[169][10]=32'h38b2e317;	data[169][11]=32'h3a0da240;	data[169][12]=32'h00000000;	data[169][13]=32'h39fd7389;	data[169][14]=32'h00000000;	data[169][15]=32'h37ee3c89;	data[169][16]=32'h38ee87b3;
data[170][0]=32'h3ade48f6;	data[170][1]=32'h3f7ffe09;	data[170][2]=32'h3bed2384;	data[170][3]=32'h00000000;	data[170][4]=32'h00000000;	data[170][5]=32'h00000000;	data[170][6]=32'h00000000;	data[170][7]=32'h00000000;	data[170][8]=32'h00000000;	data[170][9]=32'h00000000;	data[170][10]=32'h00000000;	data[170][11]=32'h00000000;	data[170][12]=32'h00000000;	data[170][13]=32'h00000000;	data[170][14]=32'h00000000;	data[170][15]=32'h00000000;	data[170][16]=32'h00000000;
data[171][0]=32'h00000000;	data[171][1]=32'h3f2baf10;	data[171][2]=32'h00000000;	data[171][3]=32'h398e7b02;	data[171][4]=32'h38fd4b45;	data[171][5]=32'h397d4b45;	data[171][6]=32'h3a2639bb;	data[171][7]=32'h387d5602;	data[171][8]=32'h00000000;	data[171][9]=32'h387d5602;	data[171][10]=32'h398e7b02;	data[171][11]=32'h38fd4b45;	data[171][12]=32'h00000000;	data[171][13]=32'h398e7b02;	data[171][14]=32'h397d4b45;	data[171][15]=32'h387d5602;	data[171][16]=32'h387d5602;
data[172][0]=32'h00000000;	data[172][1]=32'h3f1b6849;	data[172][2]=32'h00000000;	data[172][3]=32'h39b238a2;	data[172][4]=32'h00000000;	data[172][5]=32'h39819d4f;	data[172][6]=32'h38c267ef;	data[172][7]=32'h392203f6;	data[172][8]=32'h38819a9f;	data[172][9]=32'h38c267ef;	data[172][10]=32'h39b238a2;	data[172][11]=32'h00000000;	data[172][12]=32'h00000000;	data[172][13]=32'h3962d3f5;	data[172][14]=32'h39819d4f;	data[172][15]=32'h392203f6;	data[172][16]=32'h38c267ef;
data[173][0]=32'h3b3b7a95;	data[173][1]=32'h3f7ffc11;	data[173][2]=32'h3c3074a7;	data[173][3]=32'h00000000;	data[173][4]=32'h00000000;	data[173][5]=32'h390de75f;	data[173][6]=32'h00000000;	data[173][7]=32'h37e354cf;	data[173][8]=32'h00000000;	data[173][9]=32'h37e354cf;	data[173][10]=32'h00000000;	data[173][11]=32'h00000000;	data[173][12]=32'h00000000;	data[173][13]=32'h00000000;	data[173][14]=32'h390de75f;	data[173][15]=32'h37e354cf;	data[173][16]=32'h37e354cf;
data[174][0]=32'h3b43c9ef;	data[174][1]=32'h3f7ffb6a;	data[174][2]=32'h3c3c7714;	data[174][3]=32'h00000000;	data[174][4]=32'h00000000;	data[174][5]=32'h00000000;	data[174][6]=32'h38aa49eb;	data[174][7]=32'h37e354cf;	data[174][8]=32'h390de4b0;	data[174][9]=32'h37e354cf;	data[174][10]=32'h00000000;	data[174][11]=32'h00000000;	data[174][12]=32'h00000000;	data[174][13]=32'h38aa49eb;	data[174][14]=32'h00000000;	data[174][15]=32'h37e354cf;	data[174][16]=32'h37e354cf;
data[175][0]=32'h385a85f3;	data[175][1]=32'h3f205a71;	data[175][2]=32'h00000000;	data[175][3]=32'h37f4f286;	data[175][4]=32'h39c74980;	data[175][5]=32'h00000000;	data[175][6]=32'h00000000;	data[175][7]=32'h39994bec;	data[175][8]=32'h38f5486c;	data[175][9]=32'h39c74980;	data[175][10]=32'h37f4f286;	data[175][11]=32'h39c74980;	data[175][12]=32'h39b7f4f9;	data[175][13]=32'h39194d43;	data[175][14]=32'h00000000;	data[175][15]=32'h39994bec;	data[175][16]=32'h39c74980;
data[176][0]=32'h395c1df9;	data[176][1]=32'h3f1d5476;	data[176][2]=32'h00000000;	data[176][3]=32'h38b8f804;	data[176][4]=32'h3976b020;	data[176][5]=32'h38f6b020;	data[176][6]=32'h00000000;	data[176][7]=32'h39d7d970;	data[176][8]=32'h00000000;	data[176][9]=32'h00000000;	data[176][10]=32'h38b8f804;	data[176][11]=32'h3976b020;	data[176][12]=32'h00000000;	data[176][13]=32'h39c86e18;	data[176][14]=32'h38f6b020;	data[176][15]=32'h39d7d970;	data[176][16]=32'h00000000;
data[177][0]=32'h39550759;	data[177][1]=32'h3f334b73;	data[177][2]=32'h00000000;	data[177][3]=32'h3937ab28;	data[177][4]=32'h39d64821;	data[177][5]=32'h00000000;	data[177][6]=32'h00000000;	data[177][7]=32'h3874f286;	data[177][8]=32'h3874f286;	data[177][9]=32'h00000000;	data[177][10]=32'h3937ab28;	data[177][11]=32'h39d64821;	data[177][12]=32'h00000000;	data[177][13]=32'h3937ab28;	data[177][14]=32'h00000000;	data[177][15]=32'h3874f286;	data[177][16]=32'h00000000;
data[178][0]=32'h3aebd322;	data[178][1]=32'h3f7ffeb0;	data[178][2]=32'h3be25199;	data[178][3]=32'h00000000;	data[178][4]=32'h00000000;	data[178][5]=32'h00000000;	data[178][6]=32'h00000000;	data[178][7]=32'h00000000;	data[178][8]=32'h00000000;	data[178][9]=32'h00000000;	data[178][10]=32'h00000000;	data[178][11]=32'h00000000;	data[178][12]=32'h00000000;	data[178][13]=32'h00000000;	data[178][14]=32'h00000000;	data[178][15]=32'h00000000;	data[178][16]=32'h00000000;
data[179][0]=32'h3b01f538;	data[179][1]=32'h3f7ffac2;	data[179][2]=32'h3c48eac0;	data[179][3]=32'h392a6a21;	data[179][4]=32'h38aa7f9b;	data[179][5]=32'h00000000;	data[179][6]=32'h37e354cf;	data[179][7]=32'h37e354cf;	data[179][8]=32'h00000000;	data[179][9]=32'h38aa7f9b;	data[179][10]=32'h392a6a21;	data[179][11]=32'h38aa7f9b;	data[179][12]=32'h00000000;	data[179][13]=32'h37e354cf;	data[179][14]=32'h00000000;	data[179][15]=32'h37e354cf;	data[179][16]=32'h38aa7f9b;
data[180][0]=32'h385c9ed2;	data[180][1]=32'h3f1a469d;	data[180][2]=32'h00000000;	data[180][3]=32'h37f776c5;	data[180][4]=32'h39772e4a;	data[180][5]=32'h38770b65;	data[180][6]=32'h00000000;	data[180][7]=32'h38770b65;	data[180][8]=32'h00000000;	data[180][9]=32'h391a7c99;	data[180][10]=32'h37f776c5;	data[180][11]=32'h39772e4a;	data[180][12]=32'h00000000;	data[180][13]=32'h39396363;	data[180][14]=32'h38770b65;	data[180][15]=32'h38770b65;	data[180][16]=32'h391a7c99;
data[181][0]=32'h3b150abf;	data[181][1]=32'h3f7ffb6a;	data[181][2]=32'h3c386b16;	data[181][3]=32'h00000000;	data[181][4]=32'h00000000;	data[181][5]=32'h00000000;	data[181][6]=32'h00000000;	data[181][7]=32'h00000000;	data[181][8]=32'h00000000;	data[181][9]=32'h00000000;	data[181][10]=32'h00000000;	data[181][11]=32'h00000000;	data[181][12]=32'h00000000;	data[181][13]=32'h00000000;	data[181][14]=32'h00000000;	data[181][15]=32'h00000000;	data[181][16]=32'h00000000;
data[182][0]=32'h3952b8ca;	data[182][1]=32'h3f354fdf;	data[182][2]=32'h00000000;	data[182][3]=32'h00000000;	data[182][4]=32'h38f3049a;	data[182][5]=32'h37f34507;	data[182][6]=32'h00000000;	data[182][7]=32'h39a71481;	data[182][8]=32'h3988b297;	data[182][9]=32'h39c57515;	data[182][10]=32'h00000000;	data[182][11]=32'h38f3049a;	data[182][12]=32'h37f34507;	data[182][13]=32'h38f3049a;	data[182][14]=32'h37f34507;	data[182][15]=32'h39a71481;	data[182][16]=32'h39c57515;
data[183][0]=32'h00000000;	data[183][1]=32'h3f3861a6;	data[183][2]=32'h00000000;	data[183][3]=32'h00000000;	data[183][4]=32'h38f258cd;	data[183][5]=32'h39a69d0d;	data[183][6]=32'h00000000;	data[183][7]=32'h38b5d2b5;	data[183][8]=32'h00000000;	data[183][9]=32'h00000000;	data[183][10]=32'h00000000;	data[183][11]=32'h38f258cd;	data[183][12]=32'h38b5d2b5;	data[183][13]=32'h37f26e47;	data[183][14]=32'h39a69d0d;	data[183][15]=32'h38b5d2b5;	data[183][16]=32'h00000000;
data[184][0]=32'h00000000;	data[184][1]=32'h3f1a93f3;	data[184][2]=32'h00000000;	data[184][3]=32'h3876a005;	data[184][4]=32'h3976b82e;	data[184][5]=32'h00000000;	data[184][6]=32'h00000000;	data[184][7]=32'h3957e17e;	data[184][8]=32'h00000000;	data[184][9]=32'h398ac76f;	data[184][10]=32'h3876a005;	data[184][11]=32'h3976b82e;	data[184][12]=32'h37f6a005;	data[184][13]=32'h3876a005;	data[184][14]=32'h00000000;	data[184][15]=32'h3957e17e;	data[184][16]=32'h398ac76f;
data[185][0]=32'h00000000;	data[185][1]=32'h3f2736ce;	data[185][2]=32'h00000000;	data[185][3]=32'h39974c8d;	data[185][4]=32'h39b58f99;	data[185][5]=32'h00000000;	data[185][6]=32'h00000000;	data[185][7]=32'h37f26e47;	data[185][8]=32'h00000000;	data[185][9]=32'h38b59d05;	data[185][10]=32'h39974c8d;	data[185][11]=32'h39b58f99;	data[185][12]=32'h00000000;	data[185][13]=32'h38b59d05;	data[185][14]=32'h00000000;	data[185][15]=32'h37f26e47;	data[185][16]=32'h38b59d05;
data[186][0]=32'h3b136750;	data[186][1]=32'h3f7ffc11;	data[186][2]=32'h3c30079a;	data[186][3]=32'h00000000;	data[186][4]=32'h00000000;	data[186][5]=32'h00000000;	data[186][6]=32'h37e354cf;	data[186][7]=32'h00000000;	data[186][8]=32'h00000000;	data[186][9]=32'h00000000;	data[186][10]=32'h00000000;	data[186][11]=32'h00000000;	data[186][12]=32'h00000000;	data[186][13]=32'h00000000;	data[186][14]=32'h00000000;	data[186][15]=32'h00000000;	data[186][16]=32'h00000000;
data[187][0]=32'h3b1b7f4d;	data[187][1]=32'h3f7ffc11;	data[187][2]=32'h3c266dbd;	data[187][3]=32'h00000000;	data[187][4]=32'h00000000;	data[187][5]=32'h00000000;	data[187][6]=32'h00000000;	data[187][7]=32'h00000000;	data[187][8]=32'h00000000;	data[187][9]=32'h00000000;	data[187][10]=32'h00000000;	data[187][11]=32'h00000000;	data[187][12]=32'h00000000;	data[187][13]=32'h00000000;	data[187][14]=32'h00000000;	data[187][15]=32'h00000000;	data[187][16]=32'h00000000;
data[188][0]=32'h00000000;	data[188][1]=32'h3f215b57;	data[188][2]=32'h00000000;	data[188][3]=32'h00000000;	data[188][4]=32'h38798fa3;	data[188][5]=32'h38f95f52;	data[188][6]=32'h00000000;	data[188][7]=32'h00000000;	data[188][8]=32'h37f92444;	data[188][9]=32'h395a32bc;	data[188][10]=32'h00000000;	data[188][11]=32'h38798fa3;	data[188][12]=32'h391bd990;	data[188][13]=32'h38798fa3;	data[188][14]=32'h38f95f52;	data[188][15]=32'h00000000;	data[188][16]=32'h395a32bc;
data[189][0]=32'h3b542587;	data[189][1]=32'h3f7ffa1a;	data[189][2]=32'h3c4e746d;	data[189][3]=32'h00000000;	data[189][4]=32'h00000000;	data[189][5]=32'h00000000;	data[189][6]=32'h00000000;	data[189][7]=32'h00000000;	data[189][8]=32'h00000000;	data[189][9]=32'h00000000;	data[189][10]=32'h00000000;	data[189][11]=32'h00000000;	data[189][12]=32'h00000000;	data[189][13]=32'h00000000;	data[189][14]=32'h00000000;	data[189][15]=32'h00000000;	data[189][16]=32'h00000000;
data[190][0]=32'h3b296c75;	data[190][1]=32'h3f7ffcb9;	data[190][2]=32'h3c175b66;	data[190][3]=32'h00000000;	data[190][4]=32'h00000000;	data[190][5]=32'h00000000;	data[190][6]=32'h37e1a74f;	data[190][7]=32'h00000000;	data[190][8]=32'h00000000;	data[190][9]=32'h00000000;	data[190][10]=32'h00000000;	data[190][11]=32'h00000000;	data[190][12]=32'h00000000;	data[190][13]=32'h00000000;	data[190][14]=32'h00000000;	data[190][15]=32'h00000000;	data[190][16]=32'h00000000;
data[191][0]=32'h3ae56dae;	data[191][1]=32'h3f7ffeb0;	data[191][2]=32'h3bdd9572;	data[191][3]=32'h00000000;	data[191][4]=32'h00000000;	data[191][5]=32'h00000000;	data[191][6]=32'h00000000;	data[191][7]=32'h00000000;	data[191][8]=32'h00000000;	data[191][9]=32'h00000000;	data[191][10]=32'h00000000;	data[191][11]=32'h00000000;	data[191][12]=32'h00000000;	data[191][13]=32'h00000000;	data[191][14]=32'h00000000;	data[191][15]=32'h00000000;	data[191][16]=32'h00000000;
data[192][0]=32'h00000000;	data[192][1]=32'h3f1b9043;	data[192][2]=32'h00000000;	data[192][3]=32'h3878b8e4;	data[192][4]=32'h39ca0b7c;	data[192][5]=32'h00000000;	data[192][6]=32'h00000000;	data[192][7]=32'h393a7fee;	data[192][8]=32'h00000000;	data[192][9]=32'h00000000;	data[192][10]=32'h3878b8e4;	data[192][11]=32'h39ca0b7c;	data[192][12]=32'h00000000;	data[192][13]=32'h37f84d84;	data[192][14]=32'h00000000;	data[192][15]=32'h393a7fee;	data[192][16]=32'h00000000;
data[193][0]=32'h383f42a1;	data[193][1]=32'h3f2e9f6b;	data[193][2]=32'h00000000;	data[193][3]=32'h00000000;	data[193][4]=32'h00000000;	data[193][5]=32'h00000000;	data[193][6]=32'h00000000;	data[193][7]=32'h38f48c84;	data[193][8]=32'h39a82248;	data[193][9]=32'h37f4f286;	data[193][10]=32'h00000000;	data[193][11]=32'h00000000;	data[193][12]=32'h38f48c84;	data[193][13]=32'h38748726;	data[193][14]=32'h00000000;	data[193][15]=32'h38f48c84;	data[193][16]=32'h37f4f286;
data[194][0]=32'h3b211b6e;	data[194][1]=32'h3f7ffeb0;	data[194][2]=32'h3bc508b3;	data[194][3]=32'h00000000;	data[194][4]=32'h00000000;	data[194][5]=32'h37e1a74f;	data[194][6]=32'h37e1a74f;	data[194][7]=32'h00000000;	data[194][8]=32'h37e1a74f;	data[194][9]=32'h00000000;	data[194][10]=32'h00000000;	data[194][11]=32'h00000000;	data[194][12]=32'h00000000;	data[194][13]=32'h38a907cc;	data[194][14]=32'h37e1a74f;	data[194][15]=32'h00000000;	data[194][16]=32'h00000000;
data[195][0]=32'h3ac1cd95;	data[195][1]=32'h3f7ffeb0;	data[195][2]=32'h3bbb2fec;	data[195][3]=32'h00000000;	data[195][4]=32'h00000000;	data[195][5]=32'h00000000;	data[195][6]=32'h00000000;	data[195][7]=32'h00000000;	data[195][8]=32'h00000000;	data[195][9]=32'h00000000;	data[195][10]=32'h00000000;	data[195][11]=32'h00000000;	data[195][12]=32'h00000000;	data[195][13]=32'h00000000;	data[195][14]=32'h00000000;	data[195][15]=32'h00000000;	data[195][16]=32'h00000000;
data[196][0]=32'h00000000;	data[196][1]=32'h3ef0fcf8;	data[196][2]=32'h00000000;	data[196][3]=32'h00000000;	data[196][4]=32'h398ac210;	data[196][5]=32'h38b8f804;	data[196][6]=32'h00000000;	data[196][7]=32'h38b8f804;	data[196][8]=32'h38b8f804;	data[196][9]=32'h398ac210;	data[196][10]=32'h00000000;	data[196][11]=32'h398ac210;	data[196][12]=32'h398ac210;	data[196][13]=32'h38f6b020;	data[196][14]=32'h38b8f804;	data[196][15]=32'h38b8f804;	data[196][16]=32'h398ac210;
data[197][0]=32'h3b1f6083;	data[197][1]=32'h3f7ffe09;	data[197][2]=32'h3bf3519c;	data[197][3]=32'h00000000;	data[197][4]=32'h00000000;	data[197][5]=32'h00000000;	data[197][6]=32'h00000000;	data[197][7]=32'h00000000;	data[197][8]=32'h00000000;	data[197][9]=32'h00000000;	data[197][10]=32'h00000000;	data[197][11]=32'h00000000;	data[197][12]=32'h00000000;	data[197][13]=32'h00000000;	data[197][14]=32'h00000000;	data[197][15]=32'h00000000;	data[197][16]=32'h00000000;
data[198][0]=32'h38be6be1;	data[198][1]=32'h3ef692f7;	data[198][2]=32'h00000000;	data[198][3]=32'h38f5f997;	data[198][4]=32'h39a91bee;	data[198][5]=32'h3875c945;	data[198][6]=32'h37f5c945;	data[198][7]=32'h39e69a53;	data[198][8]=32'h3875c945;	data[198][9]=32'h38f5f997;	data[198][10]=32'h38f5f997;	data[198][11]=32'h39a91bee;	data[198][12]=32'h00000000;	data[198][13]=32'h39387c89;	data[198][14]=32'h3875c945;	data[198][15]=32'h39e69a53;	data[198][16]=32'h38f5f997;
data[199][0]=32'h3b126f03;	data[199][1]=32'h3f7fff58;	data[199][2]=32'h3bad71be;	data[199][3]=32'h00000000;	data[199][4]=32'h00000000;	data[199][5]=32'h00000000;	data[199][6]=32'h00000000;	data[199][7]=32'h00000000;	data[199][8]=32'h00000000;	data[199][9]=32'h00000000;	data[199][10]=32'h00000000;	data[199][11]=32'h00000000;	data[199][12]=32'h00000000;	data[199][13]=32'h00000000;	data[199][14]=32'h00000000;	data[199][15]=32'h00000000;	data[199][16]=32'h00000000;
data[200][0]=32'h00000000;	data[200][1]=32'h3f193e81;	data[200][2]=32'h00000000;	data[200][3]=32'h38cd19fa;	data[200][4]=32'h39aaf059;	data[200][5]=32'h396f5106;	data[200][6]=32'h3888bbfc;	data[200][7]=32'h3908c15a;	data[200][8]=32'h392af059;	data[200][9]=32'h39ef4faf;	data[200][10]=32'h38cd19fa;	data[200][11]=32'h39aaf059;	data[200][12]=32'h3988c003;	data[200][13]=32'h394d1f58;	data[200][14]=32'h396f5106;	data[200][15]=32'h3908c15a;	data[200][16]=32'h39ef4faf;
data[201][0]=32'h3b1aabe8;	data[201][1]=32'h3f7ffeb0;	data[201][2]=32'h3bc3cb9c;	data[201][3]=32'h00000000;	data[201][4]=32'h00000000;	data[201][5]=32'h00000000;	data[201][6]=32'h00000000;	data[201][7]=32'h00000000;	data[201][8]=32'h00000000;	data[201][9]=32'h00000000;	data[201][10]=32'h00000000;	data[201][11]=32'h00000000;	data[201][12]=32'h00000000;	data[201][13]=32'h00000000;	data[201][14]=32'h00000000;	data[201][15]=32'h00000000;	data[201][16]=32'h00000000;
data[202][0]=32'h3b25ba39;	data[202][1]=32'h3f7ffeb0;	data[202][2]=32'h3bbc91ec;	data[202][3]=32'h00000000;	data[202][4]=32'h00000000;	data[202][5]=32'h00000000;	data[202][6]=32'h00000000;	data[202][7]=32'h00000000;	data[202][8]=32'h00000000;	data[202][9]=32'h00000000;	data[202][10]=32'h00000000;	data[202][11]=32'h00000000;	data[202][12]=32'h00000000;	data[202][13]=32'h00000000;	data[202][14]=32'h00000000;	data[202][15]=32'h00000000;	data[202][16]=32'h00000000;
data[203][0]=32'h00000000;	data[203][1]=32'h3f17d0d0;	data[203][2]=32'h00000000;	data[203][3]=32'h388c825a;	data[203][4]=32'h3a41145d;	data[203][5]=32'h00000000;	data[203][6]=32'h00000000;	data[203][7]=32'h388c825a;	data[203][8]=32'h39af86c1;	data[203][9]=32'h3a41145d;	data[203][10]=32'h388c825a;	data[203][11]=32'h3a41145d;	data[203][12]=32'h39c1145d;	data[203][13]=32'h392f8818;	data[203][14]=32'h00000000;	data[203][15]=32'h388c825a;	data[203][16]=32'h3a41145d;
data[204][0]=32'h3b38a929;	data[204][1]=32'h3f7ffb6a;	data[204][2]=32'h3c3e1eb4;	data[204][3]=32'h00000000;	data[204][4]=32'h00000000;	data[204][5]=32'h00000000;	data[204][6]=32'h00000000;	data[204][7]=32'h00000000;	data[204][8]=32'h00000000;	data[204][9]=32'h00000000;	data[204][10]=32'h00000000;	data[204][11]=32'h00000000;	data[204][12]=32'h00000000;	data[204][13]=32'h00000000;	data[204][14]=32'h00000000;	data[204][15]=32'h00000000;	data[204][16]=32'h00000000;
data[205][0]=32'h00000000;	data[205][1]=32'h3f1be814;	data[205][2]=32'h00000000;	data[205][3]=32'h39b5218a;	data[205][4]=32'h39a6096a;	data[205][5]=32'h3971820e;	data[205][6]=32'h38719787;	data[205][7]=32'h3935218a;	data[205][8]=32'h00000000;	data[205][9]=32'h00000000;	data[205][10]=32'h39b5218a;	data[205][11]=32'h39a6096a;	data[205][12]=32'h37f19787;	data[205][13]=32'h39f1820e;	data[205][14]=32'h3971820e;	data[205][15]=32'h3935218a;	data[205][16]=32'h00000000;
data[206][0]=32'h3b40ab56;	data[206][1]=32'h3f7ffc11;	data[206][2]=32'h3c2d1d04;	data[206][3]=32'h386354cf;	data[206][4]=32'h392a74de;	data[206][5]=32'h38aa7f9b;	data[206][6]=32'h398e0b9c;	data[206][7]=32'h38e344b3;	data[206][8]=32'h37e354cf;	data[206][9]=32'h38e344b3;	data[206][10]=32'h386354cf;	data[206][11]=32'h392a74de;	data[206][12]=32'h386354cf;	data[206][13]=32'h39634763;	data[206][14]=32'h38aa7f9b;	data[206][15]=32'h38e344b3;	data[206][16]=32'h38e344b3;
data[207][0]=32'h3b1f6230;	data[207][1]=32'h3f7ffd61;	data[207][2]=32'h3c0feb30;	data[207][3]=32'h00000000;	data[207][4]=32'h00000000;	data[207][5]=32'h00000000;	data[207][6]=32'h00000000;	data[207][7]=32'h00000000;	data[207][8]=32'h00000000;	data[207][9]=32'h00000000;	data[207][10]=32'h00000000;	data[207][11]=32'h00000000;	data[207][12]=32'h00000000;	data[207][13]=32'h00000000;	data[207][14]=32'h00000000;	data[207][15]=32'h00000000;	data[207][16]=32'h00000000;
data[208][0]=32'h3b2181c5;	data[208][1]=32'h3f7ffcb9;	data[208][2]=32'h3c1b0b1e;	data[208][3]=32'h00000000;	data[208][4]=32'h00000000;	data[208][5]=32'h386212af;	data[208][6]=32'h37e27e0f;	data[208][7]=32'h00000000;	data[208][8]=32'h00000000;	data[208][9]=32'h00000000;	data[208][10]=32'h00000000;	data[208][11]=32'h00000000;	data[208][12]=32'h00000000;	data[208][13]=32'h37e27e0f;	data[208][14]=32'h386212af;	data[208][15]=32'h00000000;	data[208][16]=32'h00000000;
data[209][0]=32'h394125d0;	data[209][1]=32'h3f1ee243;	data[209][2]=32'h00000000;	data[209][3]=32'h38ed3ad6;	data[209][4]=32'h39de6881;	data[209][5]=32'h38b1d6a7;	data[209][6]=32'h00000000;	data[209][7]=32'h00000000;	data[209][8]=32'h00000000;	data[209][9]=32'h38ed3ad6;	data[209][10]=32'h38ed3ad6;	data[209][11]=32'h39de6881;	data[209][12]=32'h38b1d6a7;	data[209][13]=32'h3931ec21;	data[209][14]=32'h38b1d6a7;	data[209][15]=32'h00000000;	data[209][16]=32'h38ed3ad6;
data[210][0]=32'h3b2b133f;	data[210][1]=32'h3f7ffcb9;	data[210][2]=32'h3c1634f6;	data[210][3]=32'h00000000;	data[210][4]=32'h00000000;	data[210][5]=32'h00000000;	data[210][6]=32'h00000000;	data[210][7]=32'h00000000;	data[210][8]=32'h00000000;	data[210][9]=32'h00000000;	data[210][10]=32'h00000000;	data[210][11]=32'h00000000;	data[210][12]=32'h37e1a74f;	data[210][13]=32'h00000000;	data[210][14]=32'h00000000;	data[210][15]=32'h00000000;	data[210][16]=32'h00000000;
data[211][0]=32'h3b162b50;	data[211][1]=32'h3f7ffd61;	data[211][2]=32'h3c0cefd3;	data[211][3]=32'h00000000;	data[211][4]=32'h00000000;	data[211][5]=32'h00000000;	data[211][6]=32'h00000000;	data[211][7]=32'h00000000;	data[211][8]=32'h00000000;	data[211][9]=32'h00000000;	data[211][10]=32'h00000000;	data[211][11]=32'h00000000;	data[211][12]=32'h37e1a74f;	data[211][13]=32'h00000000;	data[211][14]=32'h00000000;	data[211][15]=32'h00000000;	data[211][16]=32'h00000000;
data[212][0]=32'h3946d20c;	data[212][1]=32'h3f1401a3;	data[212][2]=32'h00000000;	data[212][3]=32'h3872d9a7;	data[212][4]=32'h3a26df7d;	data[212][5]=32'h00000000;	data[212][6]=32'h00000000;	data[212][7]=32'h39a6ded2;	data[212][8]=32'h38b60865;	data[212][9]=32'h3a101dc5;	data[212][10]=32'h3872d9a7;	data[212][11]=32'h3a26df7d;	data[212][12]=32'h3a17b3e6;	data[212][13]=32'h00000000;	data[212][14]=32'h00000000;	data[212][15]=32'h39a6ded2;	data[212][16]=32'h3a101dc5;
data[213][0]=32'h3a7e67cf;	data[213][1]=32'h3f23ecab;	data[213][2]=32'h00000000;	data[213][3]=32'h39a981ef;	data[213][4]=32'h3a2981ef;	data[213][5]=32'h3876a005;	data[213][6]=32'h38b8f804;	data[213][7]=32'h3876a005;	data[213][8]=32'h00000000;	data[213][9]=32'h391a1946;	data[213][10]=32'h39a981ef;	data[213][11]=32'h3a2981ef;	data[213][12]=32'h00000000;	data[213][13]=32'h3a38eb44;	data[213][14]=32'h3876a005;	data[213][15]=32'h3876a005;	data[213][16]=32'h391a1946;
data[214][0]=32'h3ae5994c;	data[214][1]=32'h3f2396d1;	data[214][2]=32'h00000000;	data[214][3]=32'h387776c5;	data[214][4]=32'h398b4da6;	data[214][5]=32'h391ac7c2;	data[214][6]=32'h398b4da6;	data[214][7]=32'h399ac7c2;	data[214][8]=32'h3958b030;	data[214][9]=32'h387776c5;	data[214][10]=32'h387776c5;	data[214][11]=32'h398b4da6;	data[214][12]=32'h00000000;	data[214][13]=32'h39d8b187;	data[214][14]=32'h391ac7c2;	data[214][15]=32'h399ac7c2;	data[214][16]=32'h387776c5;
data[215][0]=32'h3af22475;	data[215][1]=32'h3f2f1d3f;	data[215][2]=32'h00000000;	data[215][3]=32'h3972c6dc;	data[215][4]=32'h3917bd4b;	data[215][5]=32'h00000000;	data[215][6]=32'h00000000;	data[215][7]=32'h37f26e47;	data[215][8]=32'h00000000;	data[215][9]=32'h37f26e47;	data[215][10]=32'h3972c6dc;	data[215][11]=32'h3917bd4b;	data[215][12]=32'h00000000;	data[215][13]=32'h3872d9a7;	data[215][14]=32'h00000000;	data[215][15]=32'h37f26e47;	data[215][16]=32'h37f26e47;
data[216][0]=32'h3b28ad33;	data[216][1]=32'h3f7ffb6a;	data[216][2]=32'h3c4347e9;	data[216][3]=32'h39472294;	data[216][4]=32'h37e354cf;	data[216][5]=32'h3963928c;	data[216][6]=32'h00000000;	data[216][7]=32'h392aafec;	data[216][8]=32'h37e354cf;	data[216][9]=32'h37e354cf;	data[216][10]=32'h39472294;	data[216][11]=32'h37e354cf;	data[216][12]=32'h39f1cd37;	data[216][13]=32'h38aab54b;	data[216][14]=32'h3963928c;	data[216][15]=32'h392aafec;	data[216][16]=32'h37e354cf;
data[217][0]=32'h396ef5c2;	data[217][1]=32'h3f404817;	data[217][2]=32'h00000000;	data[217][3]=32'h3950bac3;	data[217][4]=32'h39fd74e0;	data[217][5]=32'h00000000;	data[217][6]=32'h00000000;	data[217][7]=32'h00000000;	data[217][8]=32'h00000000;	data[217][9]=32'h39dfa3ea;	data[217][10]=32'h3950bac3;	data[217][11]=32'h39fd74e0;	data[217][12]=32'h37ee3c89;	data[217][13]=32'h38ee8d11;	data[217][14]=32'h00000000;	data[217][15]=32'h00000000;	data[217][16]=32'h39dfa3ea;
data[218][0]=32'h3b7ca786;	data[218][1]=32'h3f7ffa1a;	data[218][2]=32'h3c50bfa1;	data[218][3]=32'h37e42b8e;	data[218][4]=32'h37e42b8e;	data[218][5]=32'h39b9737f;	data[218][6]=32'h3980633d;	data[218][7]=32'h39643e59;	data[218][8]=32'h390ea8a5;	data[218][9]=32'h390ea8a5;	data[218][10]=32'h37e42b8e;	data[218][11]=32'h37e42b8e;	data[218][12]=32'h390ea8a5;	data[218][13]=32'h00000000;	data[218][14]=32'h39b9737f;	data[218][15]=32'h39643e59;	data[218][16]=32'h390ea8a5;
data[219][0]=32'h3afe4e4f;	data[219][1]=32'h3f7ffeb0;	data[219][2]=32'h3bc58ab9;	data[219][3]=32'h00000000;	data[219][4]=32'h00000000;	data[219][5]=32'h00000000;	data[219][6]=32'h00000000;	data[219][7]=32'h00000000;	data[219][8]=32'h00000000;	data[219][9]=32'h00000000;	data[219][10]=32'h00000000;	data[219][11]=32'h00000000;	data[219][12]=32'h00000000;	data[219][13]=32'h00000000;	data[219][14]=32'h00000000;	data[219][15]=32'h00000000;	data[219][16]=32'h00000000;
data[220][0]=32'h3b1fb10b;	data[220][1]=32'h3f7ffd61;	data[220][2]=32'h3c14954e;	data[220][3]=32'h00000000;	data[220][4]=32'h00000000;	data[220][5]=32'h00000000;	data[220][6]=32'h00000000;	data[220][7]=32'h00000000;	data[220][8]=32'h00000000;	data[220][9]=32'h00000000;	data[220][10]=32'h00000000;	data[220][11]=32'h00000000;	data[220][12]=32'h00000000;	data[220][13]=32'h00000000;	data[220][14]=32'h00000000;	data[220][15]=32'h00000000;	data[220][16]=32'h00000000;
data[221][0]=32'h3b4c8803;	data[221][1]=32'h3f7ffcb9;	data[221][2]=32'h3c21be97;	data[221][3]=32'h00000000;	data[221][4]=32'h00000000;	data[221][5]=32'h00000000;	data[221][6]=32'h00000000;	data[221][7]=32'h00000000;	data[221][8]=32'h00000000;	data[221][9]=32'h00000000;	data[221][10]=32'h00000000;	data[221][11]=32'h00000000;	data[221][12]=32'h00000000;	data[221][13]=32'h00000000;	data[221][14]=32'h00000000;	data[221][15]=32'h00000000;	data[221][16]=32'h00000000;
data[222][0]=32'h3b072cb0;	data[222][1]=32'h3f7ffe09;	data[222][2]=32'h3c00a2bd;	data[222][3]=32'h00000000;	data[222][4]=32'h00000000;	data[222][5]=32'h00000000;	data[222][6]=32'h00000000;	data[222][7]=32'h37e0d090;	data[222][8]=32'h00000000;	data[222][9]=32'h37e0d090;	data[222][10]=32'h00000000;	data[222][11]=32'h00000000;	data[222][12]=32'h00000000;	data[222][13]=32'h00000000;	data[222][14]=32'h00000000;	data[222][15]=32'h37e0d090;	data[222][16]=32'h37e0d090;
data[223][0]=32'h3ade16a1;	data[223][1]=32'h3f7fff58;	data[223][2]=32'h3b934ba2;	data[223][3]=32'h00000000;	data[223][4]=32'h00000000;	data[223][5]=32'h37dff9d0;	data[223][6]=32'h00000000;	data[223][7]=32'h00000000;	data[223][8]=32'h00000000;	data[223][9]=32'h00000000;	data[223][10]=32'h00000000;	data[223][11]=32'h00000000;	data[223][12]=32'h00000000;	data[223][13]=32'h00000000;	data[223][14]=32'h37dff9d0;	data[223][15]=32'h00000000;	data[223][16]=32'h00000000;
data[224][0]=32'h3aeea48e;	data[224][1]=32'h3f7ffe09;	data[224][2]=32'h3c01739e;	data[224][3]=32'h00000000;	data[224][4]=32'h00000000;	data[224][5]=32'h00000000;	data[224][6]=32'h00000000;	data[224][7]=32'h00000000;	data[224][8]=32'h00000000;	data[224][9]=32'h00000000;	data[224][10]=32'h00000000;	data[224][11]=32'h00000000;	data[224][12]=32'h00000000;	data[224][13]=32'h00000000;	data[224][14]=32'h00000000;	data[224][15]=32'h00000000;	data[224][16]=32'h00000000;
data[225][0]=32'h38bc88b2;	data[225][1]=32'h3f153cde;	data[225][2]=32'h00000000;	data[225][3]=32'h00000000;	data[225][4]=32'h00000000;	data[225][5]=32'h00000000;	data[225][6]=32'h00000000;	data[225][7]=32'h386c8f0a;	data[225][8]=32'h39fb859d;	data[225][9]=32'h3a2a25ae;	data[225][10]=32'h00000000;	data[225][11]=32'h00000000;	data[225][12]=32'h38b1a0f7;	data[225][13]=32'h386c8f0a;	data[225][14]=32'h00000000;	data[225][15]=32'h386c8f0a;	data[225][16]=32'h3a2a25ae;
data[226][0]=32'h3b009693;	data[226][1]=32'h3f7ffeb0;	data[226][2]=32'h3bcd4090;	data[226][3]=32'h00000000;	data[226][4]=32'h00000000;	data[226][5]=32'h00000000;	data[226][6]=32'h00000000;	data[226][7]=32'h00000000;	data[226][8]=32'h00000000;	data[226][9]=32'h00000000;	data[226][10]=32'h00000000;	data[226][11]=32'h00000000;	data[226][12]=32'h00000000;	data[226][13]=32'h00000000;	data[226][14]=32'h00000000;	data[226][15]=32'h00000000;	data[226][16]=32'h00000000;
data[227][0]=32'h3af0cad9;	data[227][1]=32'h3f7fff58;	data[227][2]=32'h3bb223d4;	data[227][3]=32'h00000000;	data[227][4]=32'h00000000;	data[227][5]=32'h00000000;	data[227][6]=32'h00000000;	data[227][7]=32'h00000000;	data[227][8]=32'h00000000;	data[227][9]=32'h00000000;	data[227][10]=32'h00000000;	data[227][11]=32'h00000000;	data[227][12]=32'h00000000;	data[227][13]=32'h00000000;	data[227][14]=32'h00000000;	data[227][15]=32'h00000000;	data[227][16]=32'h00000000;
data[228][0]=32'h3af0f31d;	data[228][1]=32'h3f7ffeb0;	data[228][2]=32'h3bbbcda1;	data[228][3]=32'h00000000;	data[228][4]=32'h00000000;	data[228][5]=32'h00000000;	data[228][6]=32'h00000000;	data[228][7]=32'h00000000;	data[228][8]=32'h00000000;	data[228][9]=32'h00000000;	data[228][10]=32'h00000000;	data[228][11]=32'h00000000;	data[228][12]=32'h00000000;	data[228][13]=32'h00000000;	data[228][14]=32'h00000000;	data[228][15]=32'h00000000;	data[228][16]=32'h00000000;
data[229][0]=32'h3acdd286;	data[229][1]=32'h3f7fff58;	data[229][2]=32'h3ba89332;	data[229][3]=32'h00000000;	data[229][4]=32'h00000000;	data[229][5]=32'h00000000;	data[229][6]=32'h00000000;	data[229][7]=32'h00000000;	data[229][8]=32'h00000000;	data[229][9]=32'h00000000;	data[229][10]=32'h00000000;	data[229][11]=32'h00000000;	data[229][12]=32'h00000000;	data[229][13]=32'h00000000;	data[229][14]=32'h00000000;	data[229][15]=32'h00000000;	data[229][16]=32'h00000000;
data[230][0]=32'h3ae789e7;	data[230][1]=32'h3f7ffeb0;	data[230][2]=32'h3bd39a46;	data[230][3]=32'h00000000;	data[230][4]=32'h00000000;	data[230][5]=32'h00000000;	data[230][6]=32'h00000000;	data[230][7]=32'h00000000;	data[230][8]=32'h00000000;	data[230][9]=32'h00000000;	data[230][10]=32'h00000000;	data[230][11]=32'h00000000;	data[230][12]=32'h00000000;	data[230][13]=32'h00000000;	data[230][14]=32'h00000000;	data[230][15]=32'h00000000;	data[230][16]=32'h00000000;
data[231][0]=32'h3b021f2a;	data[231][1]=32'h3f7ffe09;	data[231][2]=32'h3be9ee46;	data[231][3]=32'h00000000;	data[231][4]=32'h00000000;	data[231][5]=32'h00000000;	data[231][6]=32'h00000000;	data[231][7]=32'h00000000;	data[231][8]=32'h00000000;	data[231][9]=32'h00000000;	data[231][10]=32'h00000000;	data[231][11]=32'h00000000;	data[231][12]=32'h00000000;	data[231][13]=32'h00000000;	data[231][14]=32'h00000000;	data[231][15]=32'h00000000;	data[231][16]=32'h00000000;
data[232][0]=32'h3ad77ed7;	data[232][1]=32'h3f7fff58;	data[232][2]=32'h3bb2eb7a;	data[232][3]=32'h00000000;	data[232][4]=32'h00000000;	data[232][5]=32'h00000000;	data[232][6]=32'h00000000;	data[232][7]=32'h00000000;	data[232][8]=32'h00000000;	data[232][9]=32'h00000000;	data[232][10]=32'h00000000;	data[232][11]=32'h00000000;	data[232][12]=32'h00000000;	data[232][13]=32'h00000000;	data[232][14]=32'h00000000;	data[232][15]=32'h00000000;	data[232][16]=32'h00000000;
data[233][0]=32'h3ad448c2;	data[233][1]=32'h3f7ffeb0;	data[233][2]=32'h3bbc7ea1;	data[233][3]=32'h00000000;	data[233][4]=32'h00000000;	data[233][5]=32'h00000000;	data[233][6]=32'h00000000;	data[233][7]=32'h00000000;	data[233][8]=32'h00000000;	data[233][9]=32'h00000000;	data[233][10]=32'h00000000;	data[233][11]=32'h00000000;	data[233][12]=32'h00000000;	data[233][13]=32'h00000000;	data[233][14]=32'h00000000;	data[233][15]=32'h00000000;	data[233][16]=32'h00000000;
data[234][0]=32'h00000000;	data[234][1]=32'h3f296335;	data[234][2]=32'h00000000;	data[234][3]=32'h00000000;	data[234][4]=32'h00000000;	data[234][5]=32'h38b2e317;	data[234][6]=32'h3950c2d1;	data[234][7]=32'h39151e35;	data[234][8]=32'h38b2e317;	data[234][9]=32'h00000000;	data[234][10]=32'h00000000;	data[234][11]=32'h00000000;	data[234][12]=32'h00000000;	data[234][13]=32'h39951e35;	data[234][14]=32'h38b2e317;	data[234][15]=32'h39151e35;	data[234][16]=32'h00000000;
data[235][0]=32'h00000000;	data[235][1]=32'h3f34f030;	data[235][2]=32'h00000000;	data[235][3]=32'h00000000;	data[235][4]=32'h00000000;	data[235][5]=32'h38e9645d;	data[235][6]=32'h00000000;	data[235][7]=32'h00000000;	data[235][8]=32'h00000000;	data[235][9]=32'h3869340c;	data[235][10]=32'h00000000;	data[235][11]=32'h00000000;	data[235][12]=32'h00000000;	data[235][13]=32'h3911de0e;	data[235][14]=32'h38e9645d;	data[235][15]=32'h00000000;	data[235][16]=32'h3869340c;
data[236][0]=32'h3b42b51c;	data[236][1]=32'h3f7ffd61;	data[236][2]=32'h3c121f52;	data[236][3]=32'h00000000;	data[236][4]=32'h00000000;	data[236][5]=32'h00000000;	data[236][6]=32'h00000000;	data[236][7]=32'h00000000;	data[236][8]=32'h00000000;	data[236][9]=32'h00000000;	data[236][10]=32'h00000000;	data[236][11]=32'h00000000;	data[236][12]=32'h00000000;	data[236][13]=32'h00000000;	data[236][14]=32'h00000000;	data[236][15]=32'h00000000;	data[236][16]=32'h00000000;
data[237][0]=32'h383c5302;	data[237][1]=32'h3f12c7b9;	data[237][2]=32'h00000000;	data[237][3]=32'h38b2ad67;	data[237][4]=32'h00000000;	data[237][5]=32'h00000000;	data[237][6]=32'h00000000;	data[237][7]=32'h00000000;	data[237][8]=32'h00000000;	data[237][9]=32'h3914ddc8;	data[237][10]=32'h38b2ad67;	data[237][11]=32'h00000000;	data[237][12]=32'h00000000;	data[237][13]=32'h3932a559;	data[237][14]=32'h00000000;	data[237][15]=32'h00000000;	data[237][16]=32'h3914ddc8;
data[238][0]=32'h3b043d11;	data[238][1]=32'h3f7ffeb0;	data[238][2]=32'h3bd4009e;	data[238][3]=32'h00000000;	data[238][4]=32'h00000000;	data[238][5]=32'h00000000;	data[238][6]=32'h00000000;	data[238][7]=32'h00000000;	data[238][8]=32'h00000000;	data[238][9]=32'h00000000;	data[238][10]=32'h00000000;	data[238][11]=32'h00000000;	data[238][12]=32'h00000000;	data[238][13]=32'h00000000;	data[238][14]=32'h00000000;	data[238][15]=32'h00000000;	data[238][16]=32'h00000000;
data[239][0]=32'h3b1f83be;	data[239][1]=32'h3f7ffeb0;	data[239][2]=32'h3bbcc79c;	data[239][3]=32'h00000000;	data[239][4]=32'h00000000;	data[239][5]=32'h00000000;	data[239][6]=32'h00000000;	data[239][7]=32'h00000000;	data[239][8]=32'h00000000;	data[239][9]=32'h00000000;	data[239][10]=32'h00000000;	data[239][11]=32'h00000000;	data[239][12]=32'h00000000;	data[239][13]=32'h00000000;	data[239][14]=32'h00000000;	data[239][15]=32'h00000000;	data[239][16]=32'h00000000;
data[240][0]=32'h00000000;	data[240][1]=32'h3f153847;	data[240][2]=32'h3b071385;	data[240][3]=32'h3872d9a7;	data[240][4]=32'h00000000;	data[240][5]=32'h00000000;	data[240][6]=32'h00000000;	data[240][7]=32'h37f26e47;	data[240][8]=32'h00000000;	data[240][9]=32'h3872d9a7;	data[240][10]=32'h3872d9a7;	data[240][11]=32'h00000000;	data[240][12]=32'h00000000;	data[240][13]=32'h3954562e;	data[240][14]=32'h00000000;	data[240][15]=32'h37f26e47;	data[240][16]=32'h3872d9a7;
data[241][0]=32'h3b3e835e;	data[241][1]=32'h3f7ffcb9;	data[241][2]=32'h3c1bf1ce;	data[241][3]=32'h00000000;	data[241][4]=32'h00000000;	data[241][5]=32'h00000000;	data[241][6]=32'h00000000;	data[241][7]=32'h00000000;	data[241][8]=32'h00000000;	data[241][9]=32'h00000000;	data[241][10]=32'h00000000;	data[241][11]=32'h00000000;	data[241][12]=32'h00000000;	data[241][13]=32'h00000000;	data[241][14]=32'h00000000;	data[241][15]=32'h00000000;	data[241][16]=32'h00000000;
data[242][0]=32'h3b430e07;	data[242][1]=32'h3f7ffe09;	data[242][2]=32'h3bf0e17f;	data[242][3]=32'h00000000;	data[242][4]=32'h00000000;	data[242][5]=32'h00000000;	data[242][6]=32'h386212af;	data[242][7]=32'h00000000;	data[242][8]=32'h00000000;	data[242][9]=32'h00000000;	data[242][10]=32'h00000000;	data[242][11]=32'h00000000;	data[242][12]=32'h00000000;	data[242][13]=32'h00000000;	data[242][14]=32'h00000000;	data[242][15]=32'h00000000;	data[242][16]=32'h00000000;
data[243][0]=32'h3b4f652e;	data[243][1]=32'h3f7ffeb0;	data[243][2]=32'h3bde5a94;	data[243][3]=32'h00000000;	data[243][4]=32'h00000000;	data[243][5]=32'h00000000;	data[243][6]=32'h00000000;	data[243][7]=32'h00000000;	data[243][8]=32'h00000000;	data[243][9]=32'h00000000;	data[243][10]=32'h00000000;	data[243][11]=32'h00000000;	data[243][12]=32'h00000000;	data[243][13]=32'h00000000;	data[243][14]=32'h00000000;	data[243][15]=32'h00000000;	data[243][16]=32'h00000000;
data[244][0]=32'h3b516690;	data[244][1]=32'h3f7ffe09;	data[244][2]=32'h3be737b2;	data[244][3]=32'h00000000;	data[244][4]=32'h37e27e0f;	data[244][5]=32'h00000000;	data[244][6]=32'h38e23da2;	data[244][7]=32'h00000000;	data[244][8]=32'h00000000;	data[244][9]=32'h00000000;	data[244][10]=32'h00000000;	data[244][11]=32'h37e27e0f;	data[244][12]=32'h00000000;	data[244][13]=32'h00000000;	data[244][14]=32'h00000000;	data[244][15]=32'h00000000;	data[244][16]=32'h00000000;
data[245][0]=32'h3b05e07f;	data[245][1]=32'h3f7ffe09;	data[245][2]=32'h3bfe344e;	data[245][3]=32'h00000000;	data[245][4]=32'h00000000;	data[245][5]=32'h00000000;	data[245][6]=32'h00000000;	data[245][7]=32'h00000000;	data[245][8]=32'h00000000;	data[245][9]=32'h00000000;	data[245][10]=32'h00000000;	data[245][11]=32'h00000000;	data[245][12]=32'h00000000;	data[245][13]=32'h00000000;	data[245][14]=32'h00000000;	data[245][15]=32'h00000000;	data[245][16]=32'h00000000;
data[246][0]=32'h3ab516ce;	data[246][1]=32'h3f7fff58;	data[246][2]=32'h3ba3260a;	data[246][3]=32'h00000000;	data[246][4]=32'h00000000;	data[246][5]=32'h00000000;	data[246][6]=32'h00000000;	data[246][7]=32'h00000000;	data[246][8]=32'h00000000;	data[246][9]=32'h00000000;	data[246][10]=32'h00000000;	data[246][11]=32'h00000000;	data[246][12]=32'h00000000;	data[246][13]=32'h00000000;	data[246][14]=32'h00000000;	data[246][15]=32'h00000000;	data[246][16]=32'h00000000;
data[247][0]=32'h3ab1a0f7;	data[247][1]=32'h3f7fff58;	data[247][2]=32'h3b6a0acb;	data[247][3]=32'h00000000;	data[247][4]=32'h00000000;	data[247][5]=32'h00000000;	data[247][6]=32'h37dff9d0;	data[247][7]=32'h00000000;	data[247][8]=32'h00000000;	data[247][9]=32'h00000000;	data[247][10]=32'h00000000;	data[247][11]=32'h00000000;	data[247][12]=32'h00000000;	data[247][13]=32'h00000000;	data[247][14]=32'h00000000;	data[247][15]=32'h00000000;	data[247][16]=32'h00000000;
data[248][0]=32'h3a7d49ed;	data[248][1]=32'h3f800000;	data[248][2]=32'h3b2aa129;	data[248][3]=32'h00000000;	data[248][4]=32'h00000000;	data[248][5]=32'h00000000;	data[248][6]=32'h00000000;	data[248][7]=32'h00000000;	data[248][8]=32'h00000000;	data[248][9]=32'h00000000;	data[248][10]=32'h00000000;	data[248][11]=32'h00000000;	data[248][12]=32'h00000000;	data[248][13]=32'h00000000;	data[248][14]=32'h00000000;	data[248][15]=32'h00000000;	data[248][16]=32'h00000000;
data[249][0]=32'h3d04f5d3;	data[249][1]=32'h3f7faf64;	data[249][2]=32'h3c345f18;	data[249][3]=32'h39e36ba0;	data[249][4]=32'h3a179dc1;	data[249][5]=32'h3972968b;	data[249][6]=32'h38f293dc;	data[249][7]=32'h3935f03c;	data[249][8]=32'h3972968b;	data[249][9]=32'h3ad07853;	data[249][10]=32'h39e36ba0;	data[249][11]=32'h3a179dc1;	data[249][12]=32'h39b5f03c;	data[249][13]=32'h39f29533;	data[249][14]=32'h3972968b;	data[249][15]=32'h3935f03c;	data[249][16]=32'h3ad07853;
data[250][0]=32'h00000000;	data[250][1]=32'h3f44a969;	data[250][2]=32'h3bcba8e0;	data[250][3]=32'h391b3322;	data[250][4]=32'h39c9c1ab;	data[250][5]=32'h391b3322;	data[250][6]=32'h00000000;	data[250][7]=32'h39785033;	data[250][8]=32'h38ba3a23;	data[250][9]=32'h39ba3cd2;	data[250][10]=32'h391b3322;	data[250][11]=32'h39c9c1ab;	data[250][12]=32'h38ba3a23;	data[250][13]=32'h39aab7fa;	data[250][14]=32'h391b3322;	data[250][15]=32'h39785033;	data[250][16]=32'h39ba3cd2;
data[251][0]=32'h38ee41e8;	data[251][1]=32'h3ef2c27a;	data[251][2]=32'h00000000;	data[251][3]=32'h00000000;	data[251][4]=32'h00000000;	data[251][5]=32'h00000000;	data[251][6]=32'h00000000;	data[251][7]=32'h394d149b;	data[251][8]=32'h00000000;	data[251][9]=32'h386a762b;	data[251][10]=32'h00000000;	data[251][11]=32'h00000000;	data[251][12]=32'h00000000;	data[251][13]=32'h386a762b;	data[251][14]=32'h00000000;	data[251][15]=32'h394d149b;	data[251][16]=32'h386a762b;
data[252][0]=32'h3afae940;	data[252][1]=32'h3f7fff58;	data[252][2]=32'h3b9c19a7;	data[252][3]=32'h00000000;	data[252][4]=32'h00000000;	data[252][5]=32'h00000000;	data[252][6]=32'h00000000;	data[252][7]=32'h00000000;	data[252][8]=32'h00000000;	data[252][9]=32'h00000000;	data[252][10]=32'h00000000;	data[252][11]=32'h00000000;	data[252][12]=32'h00000000;	data[252][13]=32'h00000000;	data[252][14]=32'h00000000;	data[252][15]=32'h00000000;	data[252][16]=32'h00000000;
data[253][0]=32'h38e7a164;	data[253][1]=32'h3e90f909;	data[253][2]=32'h00000000;	data[253][3]=32'h00000000;	data[253][4]=32'h37eae18b;	data[253][5]=32'h00000000;	data[253][6]=32'h00000000;	data[253][7]=32'h39eab947;	data[253][8]=32'h00000000;	data[253][9]=32'h3912b4ce;	data[253][10]=32'h00000000;	data[253][11]=32'h37eae18b;	data[253][12]=32'h00000000;	data[253][13]=32'h39300ba1;	data[253][14]=32'h00000000;	data[253][15]=32'h39eab947;	data[253][16]=32'h3912b4ce;
data[254][0]=32'h3b08b8a1;	data[254][1]=32'h3f7ffeb0;	data[254][2]=32'h3bce5f74;	data[254][3]=32'h00000000;	data[254][4]=32'h00000000;	data[254][5]=32'h00000000;	data[254][6]=32'h00000000;	data[254][7]=32'h00000000;	data[254][8]=32'h00000000;	data[254][9]=32'h00000000;	data[254][10]=32'h00000000;	data[254][11]=32'h00000000;	data[254][12]=32'h00000000;	data[254][13]=32'h00000000;	data[254][14]=32'h00000000;	data[254][15]=32'h00000000;	data[254][16]=32'h00000000;
data[255][0]=32'h3adaf4ae;	data[255][1]=32'h3f7ffeb0;	data[255][2]=32'h3bb584b2;	data[255][3]=32'h00000000;	data[255][4]=32'h00000000;	data[255][5]=32'h00000000;	data[255][6]=32'h00000000;	data[255][7]=32'h00000000;	data[255][8]=32'h00000000;	data[255][9]=32'h00000000;	data[255][10]=32'h00000000;	data[255][11]=32'h00000000;	data[255][12]=32'h00000000;	data[255][13]=32'h00000000;	data[255][14]=32'h00000000;	data[255][15]=32'h00000000;	data[255][16]=32'h00000000;
data[256][0]=32'h3abb64c5;	data[256][1]=32'h3f7fff58;	data[256][2]=32'h3ba4d7bb;	data[256][3]=32'h00000000;	data[256][4]=32'h00000000;	data[256][5]=32'h00000000;	data[256][6]=32'h00000000;	data[256][7]=32'h00000000;	data[256][8]=32'h00000000;	data[256][9]=32'h00000000;	data[256][10]=32'h00000000;	data[256][11]=32'h00000000;	data[256][12]=32'h00000000;	data[256][13]=32'h00000000;	data[256][14]=32'h00000000;	data[256][15]=32'h00000000;	data[256][16]=32'h00000000;
data[257][0]=32'h383d9521;	data[257][1]=32'h3f09dc72;	data[257][2]=32'h00000000;	data[257][3]=32'h00000000;	data[257][4]=32'h37ec8f0a;	data[257][5]=32'h00000000;	data[257][6]=32'h00000000;	data[257][7]=32'h3931a0f7;	data[257][8]=32'h396cd4d5;	data[257][9]=32'h3931a0f7;	data[257][10]=32'h00000000;	data[257][11]=32'h37ec8f0a;	data[257][12]=32'h00000000;	data[257][13]=32'h3931a0f7;	data[257][14]=32'h00000000;	data[257][15]=32'h3931a0f7;	data[257][16]=32'h3931a0f7;
data[258][0]=32'h3b3fa3ef;	data[258][1]=32'h3f7ffe09;	data[258][2]=32'h3bf92012;	data[258][3]=32'h00000000;	data[258][4]=32'h00000000;	data[258][5]=32'h00000000;	data[258][6]=32'h37e1a74f;	data[258][7]=32'h00000000;	data[258][8]=32'h00000000;	data[258][9]=32'h00000000;	data[258][10]=32'h00000000;	data[258][11]=32'h00000000;	data[258][12]=32'h00000000;	data[258][13]=32'h00000000;	data[258][14]=32'h00000000;	data[258][15]=32'h00000000;	data[258][16]=32'h00000000;
data[259][0]=32'h00000000;	data[259][1]=32'h3f17a1a1;	data[259][2]=32'h00000000;	data[259][3]=32'h00000000;	data[259][4]=32'h00000000;	data[259][5]=32'h396b67c3;	data[259][6]=32'h37ebb84a;	data[259][7]=32'h3913202e;	data[259][8]=32'h38b09488;	data[259][9]=32'h38b09488;	data[259][10]=32'h00000000;	data[259][11]=32'h00000000;	data[259][12]=32'h00000000;	data[259][13]=32'h396b67c3;	data[259][14]=32'h396b67c3;	data[259][15]=32'h3913202e;	data[259][16]=32'h38b09488;
data[260][0]=32'h3b1f6739;	data[260][1]=32'h3f7ffe09;	data[260][2]=32'h3be82441;	data[260][3]=32'h00000000;	data[260][4]=32'h00000000;	data[260][5]=32'h00000000;	data[260][6]=32'h00000000;	data[260][7]=32'h00000000;	data[260][8]=32'h00000000;	data[260][9]=32'h00000000;	data[260][10]=32'h00000000;	data[260][11]=32'h00000000;	data[260][12]=32'h00000000;	data[260][13]=32'h00000000;	data[260][14]=32'h00000000;	data[260][15]=32'h00000000;	data[260][16]=32'h00000000;
data[261][0]=32'h3b1d85b7;	data[261][1]=32'h3f7ffeb0;	data[261][2]=32'h3bcb3caa;	data[261][3]=32'h00000000;	data[261][4]=32'h00000000;	data[261][5]=32'h00000000;	data[261][6]=32'h00000000;	data[261][7]=32'h00000000;	data[261][8]=32'h00000000;	data[261][9]=32'h00000000;	data[261][10]=32'h00000000;	data[261][11]=32'h00000000;	data[261][12]=32'h00000000;	data[261][13]=32'h00000000;	data[261][14]=32'h00000000;	data[261][15]=32'h00000000;	data[261][16]=32'h00000000;
data[262][0]=32'h00000000;	data[262][1]=32'h3f30bac7;	data[262][2]=32'h00000000;	data[262][3]=32'h3878b8e4;	data[262][4]=32'h39ba9c1e;	data[262][5]=32'h3a042e4d;	data[262][6]=32'h391b80fa;	data[262][7]=32'h38f8ce5d;	data[262][8]=32'h391b80fa;	data[262][9]=32'h3a2b0f38;	data[262][10]=32'h3878b8e4;	data[262][11]=32'h39ba9c1e;	data[262][12]=32'h3a3a9c1e;	data[262][13]=32'h39ca2904;	data[262][14]=32'h3a042e4d;	data[262][15]=32'h38f8ce5d;	data[262][16]=32'h3a2b0f38;
data[263][0]=32'h00000000;	data[263][1]=32'h3f3092cd;	data[263][2]=32'h00000000;	data[263][3]=32'h3a142b46;	data[263][4]=32'h39bb290b;	data[263][5]=32'h39798cf4;	data[263][6]=32'h3a42f589;	data[263][7]=32'h3a798c48;	data[263][8]=32'h39da5b00;	data[263][9]=32'h38f98a45;	data[263][10]=32'h3a142b46;	data[263][11]=32'h39bb290b;	data[263][12]=32'h38f98a45;	data[263][13]=32'h38f98a45;	data[263][14]=32'h39798cf4;	data[263][15]=32'h3a798c48;	data[263][16]=32'h38f98a45;
data[264][0]=32'h3b3b93bf;	data[264][1]=32'h3f7ffcb9;	data[264][2]=32'h3c1d741a;	data[264][3]=32'h00000000;	data[264][4]=32'h00000000;	data[264][5]=32'h392a1ef8;	data[264][6]=32'h00000000;	data[264][7]=32'h00000000;	data[264][8]=32'h00000000;	data[264][9]=32'h3862e96f;	data[264][10]=32'h00000000;	data[264][11]=32'h00000000;	data[264][12]=32'h00000000;	data[264][13]=32'h00000000;	data[264][14]=32'h392a1ef8;	data[264][15]=32'h00000000;	data[264][16]=32'h3862e96f;
data[265][0]=32'h3b05a774;	data[265][1]=32'h3f7ffe09;	data[265][2]=32'h3c049a2e;	data[265][3]=32'h00000000;	data[265][4]=32'h00000000;	data[265][5]=32'h00000000;	data[265][6]=32'h00000000;	data[265][7]=32'h00000000;	data[265][8]=32'h00000000;	data[265][9]=32'h00000000;	data[265][10]=32'h00000000;	data[265][11]=32'h00000000;	data[265][12]=32'h00000000;	data[265][13]=32'h00000000;	data[265][14]=32'h00000000;	data[265][15]=32'h00000000;	data[265][16]=32'h00000000;
data[266][0]=32'h00000000;	data[266][1]=32'h3f3a7914;	data[266][2]=32'h00000000;	data[266][3]=32'h00000000;	data[266][4]=32'h00000000;	data[266][5]=32'h37f84d84;	data[266][6]=32'h00000000;	data[266][7]=32'h3a0b96cd;	data[266][8]=32'h37f84d84;	data[266][9]=32'h00000000;	data[266][10]=32'h00000000;	data[266][11]=32'h00000000;	data[266][12]=32'h00000000;	data[266][13]=32'h00000000;	data[266][14]=32'h37f84d84;	data[266][15]=32'h3a0b96cd;	data[266][16]=32'h00000000;
data[267][0]=32'h3b3d7f52;	data[267][1]=32'h3f7ffac2;	data[267][2]=32'h3c515ad1;	data[267][3]=32'h00000000;	data[267][4]=32'h00000000;	data[267][5]=32'h00000000;	data[267][6]=32'h00000000;	data[267][7]=32'h00000000;	data[267][8]=32'h00000000;	data[267][9]=32'h00000000;	data[267][10]=32'h00000000;	data[267][11]=32'h00000000;	data[267][12]=32'h00000000;	data[267][13]=32'h00000000;	data[267][14]=32'h00000000;	data[267][15]=32'h00000000;	data[267][16]=32'h00000000;
data[268][0]=32'h00000000;	data[268][1]=32'h3f20d25f;	data[268][2]=32'h3aa8c4b0;	data[268][3]=32'h393bf50e;	data[268][4]=32'h39cb9e24;	data[268][5]=32'h00000000;	data[268][6]=32'h387a6663;	data[268][7]=32'h391ca034;	data[268][8]=32'h391ca034;	data[268][9]=32'h398cf71f;	data[268][10]=32'h393bf50e;	data[268][11]=32'h39cb9e24;	data[268][12]=32'h39fa9abb;	data[268][13]=32'h00000000;	data[268][14]=32'h00000000;	data[268][15]=32'h391ca034;	data[268][16]=32'h398cf71f;
data[269][0]=32'h3b438a2e;	data[269][1]=32'h3f7ffc11;	data[269][2]=32'h3c3a5a04;	data[269][3]=32'h00000000;	data[269][4]=32'h00000000;	data[269][5]=32'h00000000;	data[269][6]=32'h00000000;	data[269][7]=32'h00000000;	data[269][8]=32'h00000000;	data[269][9]=32'h00000000;	data[269][10]=32'h00000000;	data[269][11]=32'h00000000;	data[269][12]=32'h00000000;	data[269][13]=32'h00000000;	data[269][14]=32'h00000000;	data[269][15]=32'h00000000;	data[269][16]=32'h00000000;
data[270][0]=32'h3b4d0c8e;	data[270][1]=32'h3f7ffc11;	data[270][2]=32'h3c32b778;	data[270][3]=32'h00000000;	data[270][4]=32'h00000000;	data[270][5]=32'h00000000;	data[270][6]=32'h00000000;	data[270][7]=32'h00000000;	data[270][8]=32'h00000000;	data[270][9]=32'h00000000;	data[270][10]=32'h00000000;	data[270][11]=32'h00000000;	data[270][12]=32'h00000000;	data[270][13]=32'h00000000;	data[270][14]=32'h00000000;	data[270][15]=32'h00000000;	data[270][16]=32'h00000000;
data[271][0]=32'h3b42ba24;	data[271][1]=32'h3f7ffeb0;	data[271][2]=32'h3be3c7bb;	data[271][3]=32'h00000000;	data[271][4]=32'h00000000;	data[271][5]=32'h00000000;	data[271][6]=32'h00000000;	data[271][7]=32'h00000000;	data[271][8]=32'h00000000;	data[271][9]=32'h00000000;	data[271][10]=32'h00000000;	data[271][11]=32'h00000000;	data[271][12]=32'h00000000;	data[271][13]=32'h00000000;	data[271][14]=32'h00000000;	data[271][15]=32'h00000000;	data[271][16]=32'h00000000;
data[272][0]=32'h3b6926a0;	data[272][1]=32'h3f7ffe09;	data[272][2]=32'h3bea1e16;	data[272][3]=32'h00000000;	data[272][4]=32'h00000000;	data[272][5]=32'h00000000;	data[272][6]=32'h00000000;	data[272][7]=32'h00000000;	data[272][8]=32'h00000000;	data[272][9]=32'h00000000;	data[272][10]=32'h00000000;	data[272][11]=32'h00000000;	data[272][12]=32'h00000000;	data[272][13]=32'h00000000;	data[272][14]=32'h00000000;	data[272][15]=32'h00000000;	data[272][16]=32'h00000000;
data[273][0]=32'h3b18c3b1;	data[273][1]=32'h3f7ffeb0;	data[273][2]=32'h3bdb95bd;	data[273][3]=32'h00000000;	data[273][4]=32'h00000000;	data[273][5]=32'h00000000;	data[273][6]=32'h00000000;	data[273][7]=32'h00000000;	data[273][8]=32'h00000000;	data[273][9]=32'h00000000;	data[273][10]=32'h00000000;	data[273][11]=32'h00000000;	data[273][12]=32'h00000000;	data[273][13]=32'h00000000;	data[273][14]=32'h00000000;	data[273][15]=32'h00000000;	data[273][16]=32'h00000000;
data[274][0]=32'h3b41490b;	data[274][1]=32'h3f7ffd61;	data[274][2]=32'h3c102d75;	data[274][3]=32'h00000000;	data[274][4]=32'h00000000;	data[274][5]=32'h00000000;	data[274][6]=32'h00000000;	data[274][7]=32'h00000000;	data[274][8]=32'h00000000;	data[274][9]=32'h00000000;	data[274][10]=32'h00000000;	data[274][11]=32'h00000000;	data[274][12]=32'h00000000;	data[274][13]=32'h00000000;	data[274][14]=32'h00000000;	data[274][15]=32'h00000000;	data[274][16]=32'h00000000;
data[275][0]=32'h384308ff;	data[275][1]=32'h3f185db7;	data[275][2]=32'h3b245839;	data[275][3]=32'h00000000;	data[275][4]=32'h00000000;	data[275][5]=32'h38c3745e;	data[275][6]=32'h3802715f;	data[275][7]=32'h39c369a2;	data[275][8]=32'h3963fb3d;	data[275][9]=32'h3922d807;	data[275][10]=32'h00000000;	data[275][11]=32'h00000000;	data[275][12]=32'h00000000;	data[275][13]=32'h39c369a2;	data[275][14]=32'h38c3745e;	data[275][15]=32'h39c369a2;	data[275][16]=32'h3922d807;
data[276][0]=32'h3846cf5d;	data[276][1]=32'h3eec0ad0;	data[276][2]=32'h3b8060e3;	data[276][3]=32'h392c17a1;	data[276][4]=32'h3970ee6a;	data[276][5]=32'h388992bb;	data[276][6]=32'h00000000;	data[276][7]=32'h3a0111b8;	data[276][8]=32'h399ae29a;	data[276][9]=32'h38ce91c9;	data[276][10]=32'h392c17a1;	data[276][11]=32'h3970ee6a;	data[276][12]=32'h38ce91c9;	data[276][13]=32'h388992bb;	data[276][14]=32'h388992bb;	data[276][15]=32'h3a0111b8;	data[276][16]=32'h38ce91c9;
data[277][0]=32'h3b6fd439;	data[277][1]=32'h3f7ffd61;	data[277][2]=32'h3c09df7d;	data[277][3]=32'h00000000;	data[277][4]=32'h00000000;	data[277][5]=32'h00000000;	data[277][6]=32'h00000000;	data[277][7]=32'h00000000;	data[277][8]=32'h00000000;	data[277][9]=32'h00000000;	data[277][10]=32'h00000000;	data[277][11]=32'h00000000;	data[277][12]=32'h00000000;	data[277][13]=32'h00000000;	data[277][14]=32'h00000000;	data[277][15]=32'h00000000;	data[277][16]=32'h00000000;
data[278][0]=32'h3ae8bb40;	data[278][1]=32'h3f7ffe09;	data[278][2]=32'h3bf18d76;	data[278][3]=32'h00000000;	data[278][4]=32'h00000000;	data[278][5]=32'h00000000;	data[278][6]=32'h00000000;	data[278][7]=32'h00000000;	data[278][8]=32'h00000000;	data[278][9]=32'h00000000;	data[278][10]=32'h00000000;	data[278][11]=32'h00000000;	data[278][12]=32'h00000000;	data[278][13]=32'h00000000;	data[278][14]=32'h00000000;	data[278][15]=32'h00000000;	data[278][16]=32'h00000000;
data[279][0]=32'h3b296ac8;	data[279][1]=32'h3ee800a8;	data[279][2]=32'h00000000;	data[279][3]=32'h38048a3e;	data[279][4]=32'h39680a15;	data[279][5]=32'h39952a49;	data[279][6]=32'h398497aa;	data[279][7]=32'h3946e227;	data[279][8]=32'h39c6e37f;	data[279][9]=32'h3925bce8;	data[279][10]=32'h38048a3e;	data[279][11]=32'h39680a15;	data[279][12]=32'h38848a3e;	data[279][13]=32'h00000000;	data[279][14]=32'h39952a49;	data[279][15]=32'h3946e227;	data[279][16]=32'h3925bce8;
data[280][0]=32'h3b7d23ad;	data[280][1]=32'h3f107bdd;	data[280][2]=32'h00000000;	data[280][3]=32'h38c521de;	data[280][4]=32'h00000000;	data[280][5]=32'h3803481e;	data[280][6]=32'h00000000;	data[280][7]=32'h00000000;	data[280][8]=32'h00000000;	data[280][9]=32'h39c52f4a;	data[280][10]=32'h38c521de;	data[280][11]=32'h00000000;	data[280][12]=32'h00000000;	data[280][13]=32'h00000000;	data[280][14]=32'h3803481e;	data[280][15]=32'h00000000;	data[280][16]=32'h39c52f4a;
data[281][0]=32'h3b028226;	data[281][1]=32'h3f7ffe09;	data[281][2]=32'h3bed85aa;	data[281][3]=32'h00000000;	data[281][4]=32'h00000000;	data[281][5]=32'h00000000;	data[281][6]=32'h00000000;	data[281][7]=32'h00000000;	data[281][8]=32'h00000000;	data[281][9]=32'h00000000;	data[281][10]=32'h00000000;	data[281][11]=32'h00000000;	data[281][12]=32'h00000000;	data[281][13]=32'h00000000;	data[281][14]=32'h00000000;	data[281][15]=32'h00000000;	data[281][16]=32'h00000000;
data[282][0]=32'h3b2c76ec;	data[282][1]=32'h3efb9f56;	data[282][2]=32'h00000000;	data[282][3]=32'h39c29591;	data[282][4]=32'h3981b97e;	data[282][5]=32'h38019a9f;	data[282][6]=32'h38c29d9f;	data[282][7]=32'h39429591;	data[282][8]=32'h392226dc;	data[282][9]=32'h39e30447;	data[282][10]=32'h39c29591;	data[282][11]=32'h3981b97e;	data[282][12]=32'h3981b97e;	data[282][13]=32'h00000000;	data[282][14]=32'h38019a9f;	data[282][15]=32'h39429591;	data[282][16]=32'h39e30447;
data[283][0]=32'h3b15cf0a;	data[283][1]=32'h3f7ffd61;	data[283][2]=32'h3c1192cf;	data[283][3]=32'h00000000;	data[283][4]=32'h00000000;	data[283][5]=32'h00000000;	data[283][6]=32'h00000000;	data[283][7]=32'h00000000;	data[283][8]=32'h00000000;	data[283][9]=32'h00000000;	data[283][10]=32'h00000000;	data[283][11]=32'h00000000;	data[283][12]=32'h00000000;	data[283][13]=32'h00000000;	data[283][14]=32'h00000000;	data[283][15]=32'h00000000;	data[283][16]=32'h00000000;
data[284][0]=32'h3b3957a5;	data[284][1]=32'h3f0e238e;	data[284][2]=32'h00000000;	data[284][3]=32'h3803481e;	data[284][4]=32'h3803481e;	data[284][5]=32'h390352db;	data[284][6]=32'h38c4ec2e;	data[284][7]=32'h00000000;	data[284][8]=32'h3803481e;	data[284][9]=32'h39b49345;	data[284][10]=32'h3803481e;	data[284][11]=32'h3803481e;	data[284][12]=32'h39242a41;	data[284][13]=32'h3803481e;	data[284][14]=32'h390352db;	data[284][15]=32'h00000000;	data[284][16]=32'h39b49345;
data[285][0]=32'h3b17f1fa;	data[285][1]=32'h3f7ffd61;	data[285][2]=32'h3c068f66;	data[285][3]=32'h00000000;	data[285][4]=32'h00000000;	data[285][5]=32'h00000000;	data[285][6]=32'h00000000;	data[285][7]=32'h00000000;	data[285][8]=32'h00000000;	data[285][9]=32'h00000000;	data[285][10]=32'h00000000;	data[285][11]=32'h00000000;	data[285][12]=32'h00000000;	data[285][13]=32'h00000000;	data[285][14]=32'h00000000;	data[285][15]=32'h00000000;	data[285][16]=32'h00000000;
data[286][0]=32'h3acf4db1;	data[286][1]=32'h3f7ffe09;	data[286][2]=32'h3be419f0;	data[286][3]=32'h00000000;	data[286][4]=32'h00000000;	data[286][5]=32'h00000000;	data[286][6]=32'h00000000;	data[286][7]=32'h00000000;	data[286][8]=32'h00000000;	data[286][9]=32'h00000000;	data[286][10]=32'h00000000;	data[286][11]=32'h00000000;	data[286][12]=32'h00000000;	data[286][13]=32'h00000000;	data[286][14]=32'h00000000;	data[286][15]=32'h00000000;	data[286][16]=32'h00000000;
data[287][0]=32'h3b120c07;	data[287][1]=32'h3f7ffb6a;	data[287][2]=32'h3c309204;	data[287][3]=32'h00000000;	data[287][4]=32'h00000000;	data[287][5]=32'h00000000;	data[287][6]=32'h00000000;	data[287][7]=32'h00000000;	data[287][8]=32'h00000000;	data[287][9]=32'h00000000;	data[287][10]=32'h00000000;	data[287][11]=32'h00000000;	data[287][12]=32'h00000000;	data[287][13]=32'h00000000;	data[287][14]=32'h00000000;	data[287][15]=32'h00000000;	data[287][16]=32'h00000000;
data[288][0]=32'h3b1ef523;	data[288][1]=32'h3f7ffc11;	data[288][2]=32'h3c2dc098;	data[288][3]=32'h37e27e0f;	data[288][4]=32'h00000000;	data[288][5]=32'h00000000;	data[288][6]=32'h00000000;	data[288][7]=32'h00000000;	data[288][8]=32'h00000000;	data[288][9]=32'h00000000;	data[288][10]=32'h37e27e0f;	data[288][11]=32'h00000000;	data[288][12]=32'h00000000;	data[288][13]=32'h00000000;	data[288][14]=32'h00000000;	data[288][15]=32'h00000000;	data[288][16]=32'h00000000;
data[289][0]=32'h3acc9a78;	data[289][1]=32'h3f7ffe09;	data[289][2]=32'h3bf5fef5;	data[289][3]=32'h37e1a74f;	data[289][4]=32'h00000000;	data[289][5]=32'h00000000;	data[289][6]=32'h00000000;	data[289][7]=32'h00000000;	data[289][8]=32'h00000000;	data[289][9]=32'h00000000;	data[289][10]=32'h37e1a74f;	data[289][11]=32'h00000000;	data[289][12]=32'h00000000;	data[289][13]=32'h00000000;	data[289][14]=32'h00000000;	data[289][15]=32'h00000000;	data[289][16]=32'h00000000;
data[290][0]=32'h3b431818;	data[290][1]=32'h3f7ffb6a;	data[290][2]=32'h3c428f5c;	data[290][3]=32'h00000000;	data[290][4]=32'h00000000;	data[290][5]=32'h00000000;	data[290][6]=32'h37e27e0f;	data[290][7]=32'h00000000;	data[290][8]=32'h00000000;	data[290][9]=32'h00000000;	data[290][10]=32'h00000000;	data[290][11]=32'h00000000;	data[290][12]=32'h00000000;	data[290][13]=32'h00000000;	data[290][14]=32'h00000000;	data[290][15]=32'h00000000;	data[290][16]=32'h00000000;
data[291][0]=32'h39d3d555;	data[291][1]=32'h3f0ffac2;	data[291][2]=32'h00000000;	data[291][3]=32'h00000000;	data[291][4]=32'h39848e45;	data[291][5]=32'h00000000;	data[291][6]=32'h00000000;	data[291][7]=32'h38b0ca38;	data[291][8]=32'h38b0ca38;	data[291][9]=32'h3930bf7b;	data[291][10]=32'h00000000;	data[291][11]=32'h39848e45;	data[291][12]=32'h396ba82f;	data[291][13]=32'h00000000;	data[291][14]=32'h00000000;	data[291][15]=32'h38b0ca38;	data[291][16]=32'h3930bf7b;
data[292][0]=32'h39b823f3;	data[292][1]=32'h3eb3e187;	data[292][2]=32'h00000000;	data[292][3]=32'h00000000;	data[292][4]=32'h386d65ca;	data[292][5]=32'h39146d0a;	data[292][6]=32'h37ed65ca;	data[292][7]=32'h39146d0a;	data[292][8]=32'h00000000;	data[292][9]=32'h38b20c57;	data[292][10]=32'h00000000;	data[292][11]=32'h386d65ca;	data[292][12]=32'h00000000;	data[292][13]=32'h39946e62;	data[292][14]=32'h39146d0a;	data[292][15]=32'h39146d0a;	data[292][16]=32'h38b20c57;
data[293][0]=32'h3b10c331;	data[293][1]=32'h3f7ffeb0;	data[293][2]=32'h3bda1159;	data[293][3]=32'h00000000;	data[293][4]=32'h00000000;	data[293][5]=32'h00000000;	data[293][6]=32'h00000000;	data[293][7]=32'h00000000;	data[293][8]=32'h00000000;	data[293][9]=32'h00000000;	data[293][10]=32'h00000000;	data[293][11]=32'h00000000;	data[293][12]=32'h00000000;	data[293][13]=32'h00000000;	data[293][14]=32'h00000000;	data[293][15]=32'h00000000;	data[293][16]=32'h00000000;
data[294][0]=32'h3ae4b521;	data[294][1]=32'h3f7ffeb0;	data[294][2]=32'h3bcb9df9;	data[294][3]=32'h00000000;	data[294][4]=32'h00000000;	data[294][5]=32'h00000000;	data[294][6]=32'h00000000;	data[294][7]=32'h00000000;	data[294][8]=32'h00000000;	data[294][9]=32'h00000000;	data[294][10]=32'h00000000;	data[294][11]=32'h00000000;	data[294][12]=32'h00000000;	data[294][13]=32'h00000000;	data[294][14]=32'h00000000;	data[294][15]=32'h00000000;	data[294][16]=32'h00000000;
data[295][0]=32'h3b218a29;	data[295][1]=32'h3f7ffcb9;	data[295][2]=32'h3c260d45;	data[295][3]=32'h00000000;	data[295][4]=32'h00000000;	data[295][5]=32'h00000000;	data[295][6]=32'h00000000;	data[295][7]=32'h00000000;	data[295][8]=32'h00000000;	data[295][9]=32'h00000000;	data[295][10]=32'h00000000;	data[295][11]=32'h00000000;	data[295][12]=32'h00000000;	data[295][13]=32'h00000000;	data[295][14]=32'h00000000;	data[295][15]=32'h00000000;	data[295][16]=32'h00000000;
data[296][0]=32'h3b289408;	data[296][1]=32'h3f7ffb6a;	data[296][2]=32'h3c3a732e;	data[296][3]=32'h00000000;	data[296][4]=32'h00000000;	data[296][5]=32'h00000000;	data[296][6]=32'h00000000;	data[296][7]=32'h00000000;	data[296][8]=32'h00000000;	data[296][9]=32'h00000000;	data[296][10]=32'h00000000;	data[296][11]=32'h00000000;	data[296][12]=32'h00000000;	data[296][13]=32'h00000000;	data[296][14]=32'h00000000;	data[296][15]=32'h00000000;	data[296][16]=32'h00000000;
data[297][0]=32'h3b42efd4;	data[297][1]=32'h3f7ffa1a;	data[297][2]=32'h3c51cc10;	data[297][3]=32'h00000000;	data[297][4]=32'h00000000;	data[297][5]=32'h38aab54b;	data[297][6]=32'h3947380d;	data[297][7]=32'h3863c02e;	data[297][8]=32'h00000000;	data[297][9]=32'h3863c02e;	data[297][10]=32'h00000000;	data[297][11]=32'h00000000;	data[297][12]=32'h00000000;	data[297][13]=32'h3863c02e;	data[297][14]=32'h38aab54b;	data[297][15]=32'h3863c02e;	data[297][16]=32'h3863c02e;
data[298][0]=32'h3b204d12;	data[298][1]=32'h3f7ffcb9;	data[298][2]=32'h3c21cb97;	data[298][3]=32'h00000000;	data[298][4]=32'h00000000;	data[298][5]=32'h00000000;	data[298][6]=32'h37e354cf;	data[298][7]=32'h00000000;	data[298][8]=32'h00000000;	data[298][9]=32'h00000000;	data[298][10]=32'h00000000;	data[298][11]=32'h00000000;	data[298][12]=32'h00000000;	data[298][13]=32'h00000000;	data[298][14]=32'h00000000;	data[298][15]=32'h00000000;	data[298][16]=32'h00000000;
data[299][0]=32'h3b0ea54a;	data[299][1]=32'h3f7ffc11;	data[299][2]=32'h3c28c587;	data[299][3]=32'h00000000;	data[299][4]=32'h00000000;	data[299][5]=32'h00000000;	data[299][6]=32'h37e354cf;	data[299][7]=32'h00000000;	data[299][8]=32'h00000000;	data[299][9]=32'h00000000;	data[299][10]=32'h00000000;	data[299][11]=32'h00000000;	data[299][12]=32'h37e354cf;	data[299][13]=32'h00000000;	data[299][14]=32'h00000000;	data[299][15]=32'h00000000;	data[299][16]=32'h00000000;
data[300][0]=32'h3840f020;	data[300][1]=32'h3f4c0054;	data[300][2]=32'h00000000;	data[300][3]=32'h38734507;	data[300][4]=32'h38734507;	data[300][5]=32'h00000000;	data[300][6]=32'h00000000;	data[300][7]=32'h37f34507;	data[300][8]=32'h37f34507;	data[300][9]=32'h38734507;	data[300][10]=32'h38734507;	data[300][11]=32'h38734507;	data[300][12]=32'h00000000;	data[300][13]=32'h00000000;	data[300][14]=32'h00000000;	data[300][15]=32'h37f34507;	data[300][16]=32'h38734507;
data[301][0]=32'h3b4fe154;	data[301][1]=32'h3f7ff972;	data[301][2]=32'h3c5bdf8f;	data[301][3]=32'h00000000;	data[301][4]=32'h00000000;	data[301][5]=32'h00000000;	data[301][6]=32'h00000000;	data[301][7]=32'h00000000;	data[301][8]=32'h00000000;	data[301][9]=32'h00000000;	data[301][10]=32'h00000000;	data[301][11]=32'h00000000;	data[301][12]=32'h00000000;	data[301][13]=32'h00000000;	data[301][14]=32'h00000000;	data[301][15]=32'h00000000;	data[301][16]=32'h00000000;
data[302][0]=32'h384f32d9;	data[302][1]=32'h3f32f05a;	data[302][2]=32'h00000000;	data[302][3]=32'h37f5c945;	data[302][4]=32'h00000000;	data[302][5]=32'h00000000;	data[302][6]=32'h00000000;	data[302][7]=32'h3919a888;	data[302][8]=32'h00000000;	data[302][9]=32'h39386460;	data[302][10]=32'h37f5c945;	data[302][11]=32'h00000000;	data[302][12]=32'h00000000;	data[302][13]=32'h39571d89;	data[302][14]=32'h00000000;	data[302][15]=32'h3919a888;	data[302][16]=32'h39386460;
data[303][0]=32'h3b2ded0e;	data[303][1]=32'h3f7ffa1a;	data[303][2]=32'h3c5349bf;	data[303][3]=32'h00000000;	data[303][4]=32'h00000000;	data[303][5]=32'h00000000;	data[303][6]=32'h3863c02e;	data[303][7]=32'h3863c02e;	data[303][8]=32'h00000000;	data[303][9]=32'h00000000;	data[303][10]=32'h00000000;	data[303][11]=32'h00000000;	data[303][12]=32'h3863c02e;	data[303][13]=32'h37e354cf;	data[303][14]=32'h00000000;	data[303][15]=32'h3863c02e;	data[303][16]=32'h00000000;
data[304][0]=32'h3b3a1032;	data[304][1]=32'h3f7ffac2;	data[304][2]=32'h3c441dd2;	data[304][3]=32'h00000000;	data[304][4]=32'h00000000;	data[304][5]=32'h00000000;	data[304][6]=32'h00000000;	data[304][7]=32'h00000000;	data[304][8]=32'h00000000;	data[304][9]=32'h00000000;	data[304][10]=32'h00000000;	data[304][11]=32'h00000000;	data[304][12]=32'h00000000;	data[304][13]=32'h00000000;	data[304][14]=32'h00000000;	data[304][15]=32'h00000000;	data[304][16]=32'h00000000;
data[305][0]=32'h3b39742a;	data[305][1]=32'h3f7ffcb9;	data[305][2]=32'h3c24fca4;	data[305][3]=32'h00000000;	data[305][4]=32'h00000000;	data[305][5]=32'h00000000;	data[305][6]=32'h00000000;	data[305][7]=32'h00000000;	data[305][8]=32'h00000000;	data[305][9]=32'h00000000;	data[305][10]=32'h00000000;	data[305][11]=32'h00000000;	data[305][12]=32'h00000000;	data[305][13]=32'h00000000;	data[305][14]=32'h00000000;	data[305][15]=32'h00000000;	data[305][16]=32'h00000000;
data[306][0]=32'h3b27b840;	data[306][1]=32'h3f7ffd61;	data[306][2]=32'h3c16d026;	data[306][3]=32'h00000000;	data[306][4]=32'h00000000;	data[306][5]=32'h00000000;	data[306][6]=32'h00000000;	data[306][7]=32'h00000000;	data[306][8]=32'h00000000;	data[306][9]=32'h00000000;	data[306][10]=32'h00000000;	data[306][11]=32'h00000000;	data[306][12]=32'h00000000;	data[306][13]=32'h00000000;	data[306][14]=32'h00000000;	data[306][15]=32'h00000000;	data[306][16]=32'h00000000;
data[307][0]=32'h3b346349;	data[307][1]=32'h3f7ffd61;	data[307][2]=32'h3c0a11d2;	data[307][3]=32'h00000000;	data[307][4]=32'h00000000;	data[307][5]=32'h00000000;	data[307][6]=32'h00000000;	data[307][7]=32'h00000000;	data[307][8]=32'h00000000;	data[307][9]=32'h00000000;	data[307][10]=32'h00000000;	data[307][11]=32'h00000000;	data[307][12]=32'h37e1a74f;	data[307][13]=32'h00000000;	data[307][14]=32'h00000000;	data[307][15]=32'h00000000;	data[307][16]=32'h00000000;
data[308][0]=32'h3b34d70d;	data[308][1]=32'h3f7ffc11;	data[308][2]=32'h3c270d20;	data[308][3]=32'h00000000;	data[308][4]=32'h00000000;	data[308][5]=32'h00000000;	data[308][6]=32'h00000000;	data[308][7]=32'h00000000;	data[308][8]=32'h00000000;	data[308][9]=32'h00000000;	data[308][10]=32'h00000000;	data[308][11]=32'h00000000;	data[308][12]=32'h00000000;	data[308][13]=32'h00000000;	data[308][14]=32'h00000000;	data[308][15]=32'h00000000;	data[308][16]=32'h00000000;
data[309][0]=32'h3b3d18fb;	data[309][1]=32'h3f7ffb6a;	data[309][2]=32'h3c3f93ff;	data[309][3]=32'h00000000;	data[309][4]=32'h00000000;	data[309][5]=32'h00000000;	data[309][6]=32'h00000000;	data[309][7]=32'h00000000;	data[309][8]=32'h00000000;	data[309][9]=32'h00000000;	data[309][10]=32'h00000000;	data[309][11]=32'h00000000;	data[309][12]=32'h00000000;	data[309][13]=32'h00000000;	data[309][14]=32'h00000000;	data[309][15]=32'h00000000;	data[309][16]=32'h00000000;
data[310][0]=32'h00000000;	data[310][1]=32'h3f001451;	data[310][2]=32'h00000000;	data[310][3]=32'h38b63e15;	data[310][4]=32'h39549bf9;	data[310][5]=32'h00000000;	data[310][6]=32'h00000000;	data[310][7]=32'h38f2f9dd;	data[310][8]=32'h38f2f9dd;	data[310][9]=32'h38b63e15;	data[310][10]=32'h38b63e15;	data[310][11]=32'h39549bf9;	data[310][12]=32'h38b63e15;	data[310][13]=32'h3872d9a7;	data[310][14]=32'h00000000;	data[310][15]=32'h38f2f9dd;	data[310][16]=32'h38b63e15;
data[311][0]=32'h3b6fa89a;	data[311][1]=32'h3f7ffc11;	data[311][2]=32'h3c3035bd;	data[311][3]=32'h00000000;	data[311][4]=32'h3862e96f;	data[311][5]=32'h00000000;	data[311][6]=32'h00000000;	data[311][7]=32'h00000000;	data[311][8]=32'h37e354cf;	data[311][9]=32'h00000000;	data[311][10]=32'h00000000;	data[311][11]=32'h3862e96f;	data[311][12]=32'h00000000;	data[311][13]=32'h00000000;	data[311][14]=32'h00000000;	data[311][15]=32'h00000000;	data[311][16]=32'h00000000;
data[312][0]=32'h3b2e9b89;	data[312][1]=32'h3f7ffeb0;	data[312][2]=32'h3bdb4104;	data[312][3]=32'h00000000;	data[312][4]=32'h38a9de8b;	data[312][5]=32'h38627e0f;	data[312][6]=32'h37e27e0f;	data[312][7]=32'h38627e0f;	data[312][8]=32'h00000000;	data[312][9]=32'h00000000;	data[312][10]=32'h00000000;	data[312][11]=32'h38a9de8b;	data[312][12]=32'h38e278b1;	data[312][13]=32'h00000000;	data[312][14]=32'h38627e0f;	data[312][15]=32'h38627e0f;	data[312][16]=32'h00000000;
data[313][0]=32'h3b85dfa8;	data[313][1]=32'h3f7ffb6a;	data[313][2]=32'h3c38a19d;	data[313][3]=32'h390dfcd8;	data[313][4]=32'h37e354cf;	data[313][5]=32'h37e354cf;	data[313][6]=32'h37e354cf;	data[313][7]=32'h38e32f3a;	data[313][8]=32'h00000000;	data[313][9]=32'h00000000;	data[313][10]=32'h390dfcd8;	data[313][11]=32'h37e354cf;	data[313][12]=32'h00000000;	data[313][13]=32'h00000000;	data[313][14]=32'h37e354cf;	data[313][15]=32'h38e32f3a;	data[313][16]=32'h00000000;
data[314][0]=32'h3b2d70e7;	data[314][1]=32'h3f7ffc11;	data[314][2]=32'h3c195ee1;	data[314][3]=32'h00000000;	data[314][4]=32'h00000000;	data[314][5]=32'h00000000;	data[314][6]=32'h390e1252;	data[314][7]=32'h00000000;	data[314][8]=32'h00000000;	data[314][9]=32'h00000000;	data[314][10]=32'h00000000;	data[314][11]=32'h00000000;	data[314][12]=32'h00000000;	data[314][13]=32'h00000000;	data[314][14]=32'h00000000;	data[314][15]=32'h00000000;	data[314][16]=32'h00000000;
data[315][0]=32'h3b18b9a0;	data[315][1]=32'h3f7ffb6a;	data[315][2]=32'h3c2f46aa;	data[315][3]=32'h00000000;	data[315][4]=32'h00000000;	data[315][5]=32'h00000000;	data[315][6]=32'h00000000;	data[315][7]=32'h00000000;	data[315][8]=32'h00000000;	data[315][9]=32'h00000000;	data[315][10]=32'h00000000;	data[315][11]=32'h00000000;	data[315][12]=32'h00000000;	data[315][13]=32'h00000000;	data[315][14]=32'h00000000;	data[315][15]=32'h00000000;	data[315][16]=32'h00000000;
data[316][0]=32'h3b0b75ea;	data[316][1]=32'h3f7ffcb9;	data[316][2]=32'h3c105a56;	data[316][3]=32'h00000000;	data[316][4]=32'h00000000;	data[316][5]=32'h00000000;	data[316][6]=32'h00000000;	data[316][7]=32'h00000000;	data[316][8]=32'h00000000;	data[316][9]=32'h00000000;	data[316][10]=32'h00000000;	data[316][11]=32'h00000000;	data[316][12]=32'h00000000;	data[316][13]=32'h00000000;	data[316][14]=32'h00000000;	data[316][15]=32'h00000000;	data[316][16]=32'h00000000;
data[317][0]=32'h3859af33;	data[317][1]=32'h3f161a61;	data[317][2]=32'h00000000;	data[317][3]=32'h3970500a;	data[317][4]=32'h39c3415e;	data[317][5]=32'h00000000;	data[317][6]=32'h00000000;	data[317][7]=32'h00000000;	data[317][8]=32'h00000000;	data[317][9]=32'h391632b2;	data[317][10]=32'h3970500a;	data[317][11]=32'h39c3415e;	data[317][12]=32'h00000000;	data[317][13]=32'h39872d5b;	data[317][14]=32'h00000000;	data[317][15]=32'h00000000;	data[317][16]=32'h391632b2;
data[318][0]=32'h39461e32;	data[318][1]=32'h3f0fd36f;	data[318][2]=32'h00000000;	data[318][3]=32'h39a06d48;	data[318][4]=32'h39e09988;	data[318][5]=32'h38805880;	data[318][6]=32'h39005880;	data[318][7]=32'h00000000;	data[318][8]=32'h00000000;	data[318][9]=32'h3a18686c;	data[318][10]=32'h39a06d48;	data[318][11]=32'h39e09988;	data[318][12]=32'h3a28737c;	data[318][13]=32'h39b07858;	data[318][14]=32'h38805880;	data[318][15]=32'h00000000;	data[318][16]=32'h3a18686c;
data[319][0]=32'h3af959f4;	data[319][1]=32'h3f7ffd61;	data[319][2]=32'h3c173033;	data[319][3]=32'h00000000;	data[319][4]=32'h00000000;	data[319][5]=32'h00000000;	data[319][6]=32'h00000000;	data[319][7]=32'h00000000;	data[319][8]=32'h00000000;	data[319][9]=32'h00000000;	data[319][10]=32'h00000000;	data[319][11]=32'h00000000;	data[319][12]=32'h00000000;	data[319][13]=32'h00000000;	data[319][14]=32'h00000000;	data[319][15]=32'h00000000;	data[319][16]=32'h00000000;
data[320][0]=32'h3af2e713;	data[320][1]=32'h3f7ffcb9;	data[320][2]=32'h3c1f31f4;	data[320][3]=32'h00000000;	data[320][4]=32'h00000000;	data[320][5]=32'h00000000;	data[320][6]=32'h00000000;	data[320][7]=32'h00000000;	data[320][8]=32'h00000000;	data[320][9]=32'h00000000;	data[320][10]=32'h00000000;	data[320][11]=32'h00000000;	data[320][12]=32'h00000000;	data[320][13]=32'h00000000;	data[320][14]=32'h00000000;	data[320][15]=32'h00000000;	data[320][16]=32'h00000000;
data[321][0]=32'h39de8cbe;	data[321][1]=32'h3f16c02f;	data[321][2]=32'h00000000;	data[321][3]=32'h00000000;	data[321][4]=32'h00000000;	data[321][5]=32'h39bc194b;	data[321][6]=32'h38bc1d52;	data[321][7]=32'h393c17f4;	data[321][8]=32'h399cbf13;	data[321][9]=32'h395b722c;	data[321][10]=32'h00000000;	data[321][11]=32'h00000000;	data[321][12]=32'h398d11f7;	data[321][13]=32'h39ac6c2f;	data[321][14]=32'h39bc194b;	data[321][15]=32'h393c17f4;	data[321][16]=32'h395b722c;
data[322][0]=32'h3973c082;	data[322][1]=32'h3f2e4064;	data[322][2]=32'h00000000;	data[322][3]=32'h3978685c;	data[322][4]=32'h39e8e384;	data[322][5]=32'h00000000;	data[322][6]=32'h00000000;	data[322][7]=32'h00000000;	data[322][8]=32'h38784d84;	data[322][9]=32'h3a2304fd;	data[322][10]=32'h3978685c;	data[322][11]=32'h39e8e384;	data[322][12]=32'h3a49d5cc;	data[322][13]=32'h38ba3a23;	data[322][14]=32'h00000000;	data[322][15]=32'h00000000;	data[322][16]=32'h3a2304fd;
data[323][0]=32'h39c4c13b;	data[323][1]=32'h3f125c3e;	data[323][2]=32'h00000000;	data[323][3]=32'h3a269bb6;	data[323][4]=32'h39fde198;	data[323][5]=32'h00000000;	data[323][6]=32'h00000000;	data[323][7]=32'h00000000;	data[323][8]=32'h395e240d;	data[323][9]=32'h399eacff;	data[323][10]=32'h3a269bb6;	data[323][11]=32'h39fde198;	data[323][12]=32'h39fde198;	data[323][13]=32'h39fde198;	data[323][14]=32'h00000000;	data[323][15]=32'h00000000;	data[323][16]=32'h399eacff;
data[324][0]=32'h3b3dac9e;	data[324][1]=32'h3f7ffac2;	data[324][2]=32'h3c539da1;	data[324][3]=32'h00000000;	data[324][4]=32'h00000000;	data[324][5]=32'h00000000;	data[324][6]=32'h00000000;	data[324][7]=32'h00000000;	data[324][8]=32'h00000000;	data[324][9]=32'h00000000;	data[324][10]=32'h00000000;	data[324][11]=32'h00000000;	data[324][12]=32'h00000000;	data[324][13]=32'h00000000;	data[324][14]=32'h00000000;	data[324][15]=32'h00000000;	data[324][16]=32'h00000000;
data[325][0]=32'h3b0a6117;	data[325][1]=32'h3f7ffeb0;	data[325][2]=32'h3bc9cd3e;	data[325][3]=32'h00000000;	data[325][4]=32'h00000000;	data[325][5]=32'h00000000;	data[325][6]=32'h00000000;	data[325][7]=32'h00000000;	data[325][8]=32'h00000000;	data[325][9]=32'h00000000;	data[325][10]=32'h00000000;	data[325][11]=32'h00000000;	data[325][12]=32'h00000000;	data[325][13]=32'h00000000;	data[325][14]=32'h00000000;	data[325][15]=32'h00000000;	data[325][16]=32'h00000000;
data[326][0]=32'h3ac7f349;	data[326][1]=32'h3f7fff58;	data[326][2]=32'h3ba8170b;	data[326][3]=32'h00000000;	data[326][4]=32'h00000000;	data[326][5]=32'h00000000;	data[326][6]=32'h00000000;	data[326][7]=32'h00000000;	data[326][8]=32'h00000000;	data[326][9]=32'h00000000;	data[326][10]=32'h00000000;	data[326][11]=32'h00000000;	data[326][12]=32'h00000000;	data[326][13]=32'h00000000;	data[326][14]=32'h00000000;	data[326][15]=32'h00000000;	data[326][16]=32'h00000000;
data[327][0]=32'h3b9c23b8;	data[327][1]=32'h3f7ffac2;	data[327][2]=32'h3c21fa26;	data[327][3]=32'h00000000;	data[327][4]=32'h39815e39;	data[327][5]=32'h38ac987a;	data[327][6]=32'h00000000;	data[327][7]=32'h3865d90d;	data[327][8]=32'h3865d90d;	data[327][9]=32'h3865d90d;	data[327][10]=32'h00000000;	data[327][11]=32'h39815e39;	data[327][12]=32'h00000000;	data[327][13]=32'h00000000;	data[327][14]=32'h38ac987a;	data[327][15]=32'h3865d90d;	data[327][16]=32'h3865d90d;
data[328][0]=32'h00000000;	data[328][1]=32'h3f11ceaf;	data[328][2]=32'h00000000;	data[328][3]=32'h38705568;	data[328][4]=32'h38b45ae6;	data[328][5]=32'h39525827;	data[328][6]=32'h00000000;	data[328][7]=32'h39ff6c31;	data[328][8]=32'h38f06583;	data[328][9]=32'h39873970;	data[328][10]=32'h38705568;	data[328][11]=32'h38b45ae6;	data[328][12]=32'h00000000;	data[328][13]=32'h39344acb;	data[328][14]=32'h39525827;	data[328][15]=32'h39ff6c31;	data[328][16]=32'h39873970;
data[329][0]=32'h3ba623ec;	data[329][1]=32'h3f7ffa1a;	data[329][2]=32'h3c3a40d9;	data[329][3]=32'h00000000;	data[329][4]=32'h00000000;	data[329][5]=32'h00000000;	data[329][6]=32'h39650fba;	data[329][7]=32'h392bc9c8;	data[329][8]=32'h00000000;	data[329][9]=32'h00000000;	data[329][10]=32'h00000000;	data[329][11]=32'h00000000;	data[329][12]=32'h00000000;	data[329][13]=32'h37e5024e;	data[329][14]=32'h00000000;	data[329][15]=32'h392bc9c8;	data[329][16]=32'h00000000;
data[330][0]=32'h00000000;	data[330][1]=32'h3f0a1b5c;	data[330][2]=32'h00000000;	data[330][3]=32'h38b4c646;	data[330][4]=32'h39a5a76f;	data[330][5]=32'h3970f3c9;	data[330][6]=32'h3870c0c8;	data[330][7]=32'h39a5a76f;	data[330][8]=32'h3970f3c9;	data[330][9]=32'h391698b3;	data[330][10]=32'h38b4c646;	data[330][11]=32'h39a5a76f;	data[330][12]=32'h00000000;	data[330][13]=32'h39f0f3c9;	data[330][14]=32'h3970f3c9;	data[330][15]=32'h39a5a76f;	data[330][16]=32'h391698b3;
data[331][0]=32'h3b66ce00;	data[331][1]=32'h3f7ffcb9;	data[331][2]=32'h3c0df8e7;	data[331][3]=32'h37e42b8e;	data[331][4]=32'h37e42b8e;	data[331][5]=32'h38e4669c;	data[331][6]=32'h37e42b8e;	data[331][7]=32'h00000000;	data[331][8]=32'h00000000;	data[331][9]=32'h00000000;	data[331][10]=32'h37e42b8e;	data[331][11]=32'h37e42b8e;	data[331][12]=32'h00000000;	data[331][13]=32'h386496ee;	data[331][14]=32'h38e4669c;	data[331][15]=32'h00000000;	data[331][16]=32'h00000000;
data[332][0]=32'h3bcb60bc;	data[332][1]=32'h3f7ffa1a;	data[332][2]=32'h3c2c9f30;	data[332][3]=32'h00000000;	data[332][4]=32'h399e3184;	data[332][5]=32'h37e5d90d;	data[332][6]=32'h38e6197a;	data[332][7]=32'h3966197a;	data[332][8]=32'h00000000;	data[332][9]=32'h390fcfec;	data[332][10]=32'h00000000;	data[332][11]=32'h399e3184;	data[332][12]=32'h38ac987a;	data[332][13]=32'h00000000;	data[332][14]=32'h37e5d90d;	data[332][15]=32'h3966197a;	data[332][16]=32'h390fcfec;
data[333][0]=32'h3b68518e;	data[333][1]=32'h3f7ffcb9;	data[333][2]=32'h3c176f1d;	data[333][3]=32'h00000000;	data[333][4]=32'h00000000;	data[333][5]=32'h00000000;	data[333][6]=32'h38642b8e;	data[333][7]=32'h37e42b8e;	data[333][8]=32'h00000000;	data[333][9]=32'h37e42b8e;	data[333][10]=32'h00000000;	data[333][11]=32'h00000000;	data[333][12]=32'h00000000;	data[333][13]=32'h00000000;	data[333][14]=32'h00000000;	data[333][15]=32'h37e42b8e;	data[333][16]=32'h37e42b8e;
data[334][0]=32'h00000000;	data[334][1]=32'h3f0cfd4c;	data[334][2]=32'h00000000;	data[334][3]=32'h39e191d6;	data[334][4]=32'h399661ac;	data[334][5]=32'h00000000;	data[334][6]=32'h00000000;	data[334][7]=32'h39c37f1b;	data[334][8]=32'h00000000;	data[334][9]=32'h38f09b33;	data[334][10]=32'h39e191d6;	data[334][11]=32'h399661ac;	data[334][12]=32'h38b45ae6;	data[334][13]=32'h39528879;	data[334][14]=32'h00000000;	data[334][15]=32'h39c37f1b;	data[334][16]=32'h38f09b33;
data[335][0]=32'h397de447;	data[335][1]=32'h3f11bef5;	data[335][2]=32'h00000000;	data[335][3]=32'h00000000;	data[335][4]=32'h00000000;	data[335][5]=32'h38b88ca4;	data[335][6]=32'h00000000;	data[335][7]=32'h39e68f97;	data[335][8]=32'h393871cc;	data[335][9]=32'h3919b5f4;	data[335][10]=32'h00000000;	data[335][11]=32'h00000000;	data[335][12]=32'h00000000;	data[335][13]=32'h39b87324;	data[335][14]=32'h38b88ca4;	data[335][15]=32'h39e68f97;	data[335][16]=32'h3919b5f4;
data[336][0]=32'h3b1fef1e;	data[336][1]=32'h3f7ffd61;	data[336][2]=32'h3c135c69;	data[336][3]=32'h00000000;	data[336][4]=32'h386212af;	data[336][5]=32'h00000000;	data[336][6]=32'h00000000;	data[336][7]=32'h00000000;	data[336][8]=32'h00000000;	data[336][9]=32'h386212af;	data[336][10]=32'h00000000;	data[336][11]=32'h386212af;	data[336][12]=32'h00000000;	data[336][13]=32'h00000000;	data[336][14]=32'h00000000;	data[336][15]=32'h00000000;	data[336][16]=32'h386212af;
data[337][0]=32'h3b219c9d;	data[337][1]=32'h3f7ffcb9;	data[337][2]=32'h3c17c07c;	data[337][3]=32'h00000000;	data[337][4]=32'h3929f405;	data[337][5]=32'h00000000;	data[337][6]=32'h390da194;	data[337][7]=32'h00000000;	data[337][8]=32'h38627e0f;	data[337][9]=32'h37e27e0f;	data[337][10]=32'h00000000;	data[337][11]=32'h3929f405;	data[337][12]=32'h00000000;	data[337][13]=32'h37e27e0f;	data[337][14]=32'h00000000;	data[337][15]=32'h00000000;	data[337][16]=32'h37e27e0f;
data[338][0]=32'h3918fcbc;	data[338][1]=32'h3f07f8cb;	data[338][2]=32'h00000000;	data[338][3]=32'h391cd335;	data[338][4]=32'h00000000;	data[338][5]=32'h37fad1c3;	data[338][6]=32'h37fad1c3;	data[338][7]=32'h398d236a;	data[338][8]=32'h37fad1c3;	data[338][9]=32'h391cd335;	data[338][10]=32'h391cd335;	data[338][11]=32'h00000000;	data[338][12]=32'h00000000;	data[338][13]=32'h393c301c;	data[338][14]=32'h37fad1c3;	data[338][15]=32'h398d236a;	data[338][16]=32'h391cd335;
data[339][0]=32'h3b027815;	data[339][1]=32'h3f7ffeb0;	data[339][2]=32'h3bdcd482;	data[339][3]=32'h00000000;	data[339][4]=32'h00000000;	data[339][5]=32'h00000000;	data[339][6]=32'h00000000;	data[339][7]=32'h00000000;	data[339][8]=32'h00000000;	data[339][9]=32'h00000000;	data[339][10]=32'h00000000;	data[339][11]=32'h00000000;	data[339][12]=32'h00000000;	data[339][13]=32'h00000000;	data[339][14]=32'h00000000;	data[339][15]=32'h00000000;	data[339][16]=32'h00000000;
data[340][0]=32'h3ae1ae05;	data[340][1]=32'h3f7ffeb0;	data[340][2]=32'h3bd002e2;	data[340][3]=32'h00000000;	data[340][4]=32'h00000000;	data[340][5]=32'h00000000;	data[340][6]=32'h00000000;	data[340][7]=32'h00000000;	data[340][8]=32'h00000000;	data[340][9]=32'h00000000;	data[340][10]=32'h00000000;	data[340][11]=32'h00000000;	data[340][12]=32'h00000000;	data[340][13]=32'h00000000;	data[340][14]=32'h00000000;	data[340][15]=32'h00000000;	data[340][16]=32'h00000000;
data[341][0]=32'h3b3385d4;	data[341][1]=32'h3f7ffc11;	data[341][2]=32'h3c2d7d7c;	data[341][3]=32'h00000000;	data[341][4]=32'h38aa49eb;	data[341][5]=32'h37e354cf;	data[341][6]=32'h392a3c7f;	data[341][7]=32'h00000000;	data[341][8]=32'h3862e96f;	data[341][9]=32'h37e354cf;	data[341][10]=32'h00000000;	data[341][11]=32'h38aa49eb;	data[341][12]=32'h00000000;	data[341][13]=32'h00000000;	data[341][14]=32'h37e354cf;	data[341][15]=32'h00000000;	data[341][16]=32'h37e354cf;
data[342][0]=32'h3b0d9077;	data[342][1]=32'h3f7ffeb0;	data[342][2]=32'h3bccc972;	data[342][3]=32'h00000000;	data[342][4]=32'h00000000;	data[342][5]=32'h00000000;	data[342][6]=32'h37e0d090;	data[342][7]=32'h00000000;	data[342][8]=32'h00000000;	data[342][9]=32'h00000000;	data[342][10]=32'h00000000;	data[342][11]=32'h00000000;	data[342][12]=32'h00000000;	data[342][13]=32'h00000000;	data[342][14]=32'h00000000;	data[342][15]=32'h00000000;	data[342][16]=32'h00000000;
data[343][0]=32'h3849539c;	data[343][1]=32'h3f1a0f91;	data[343][2]=32'h00000000;	data[343][3]=32'h38770b65;	data[343][4]=32'h38b96363;	data[343][5]=32'h00000000;	data[343][6]=32'h00000000;	data[343][7]=32'h00000000;	data[343][8]=32'h00000000;	data[343][9]=32'h38f720de;	data[343][10]=32'h38770b65;	data[343][11]=32'h38b96363;	data[343][12]=32'h393958a7;	data[343][13]=32'h391a748b;	data[343][14]=32'h00000000;	data[343][15]=32'h00000000;	data[343][16]=32'h38f720de;
data[344][0]=32'h3b36da1c;	data[344][1]=32'h3f7ffa1a;	data[344][2]=32'h3c5b2b34;	data[344][3]=32'h00000000;	data[344][4]=32'h37e27e0f;	data[344][5]=32'h00000000;	data[344][6]=32'h397f0381;	data[344][7]=32'h37e27e0f;	data[344][8]=32'h00000000;	data[344][9]=32'h00000000;	data[344][10]=32'h00000000;	data[344][11]=32'h37e27e0f;	data[344][12]=32'h00000000;	data[344][13]=32'h00000000;	data[344][14]=32'h00000000;	data[344][15]=32'h37e27e0f;	data[344][16]=32'h00000000;
data[345][0]=32'h3b1ac00a;	data[345][1]=32'h3f7ffcb9;	data[345][2]=32'h3c1addd2;	data[345][3]=32'h00000000;	data[345][4]=32'h37e0d090;	data[345][5]=32'h00000000;	data[345][6]=32'h00000000;	data[345][7]=32'h00000000;	data[345][8]=32'h38613bf0;	data[345][9]=32'h00000000;	data[345][10]=32'h00000000;	data[345][11]=32'h37e0d090;	data[345][12]=32'h00000000;	data[345][13]=32'h00000000;	data[345][14]=32'h00000000;	data[345][15]=32'h00000000;	data[345][16]=32'h00000000;
data[346][0]=32'h3ab520df;	data[346][1]=32'h3ecdee78;	data[346][2]=32'h00000000;	data[346][3]=32'h37fe2cc1;	data[346][4]=32'h397e6271;	data[346][5]=32'h00000000;	data[346][6]=32'h37fe2cc1;	data[346][7]=32'h399efc2f;	data[346][8]=32'h00000000;	data[346][9]=32'h39ceaf50;	data[346][10]=32'h37fe2cc1;	data[346][11]=32'h397e6271;	data[346][12]=32'h393ec9d5;	data[346][13]=32'h38bed741;	data[346][14]=32'h00000000;	data[346][15]=32'h399efc2f;	data[346][16]=32'h39ceaf50;
data[347][0]=32'h00000000;	data[347][1]=32'h3f178c00;	data[347][2]=32'h00000000;	data[347][3]=32'h38f7d209;	data[347][4]=32'h39aa60bc;	data[347][5]=32'h00000000;	data[347][6]=32'h00000000;	data[347][7]=32'h00000000;	data[347][8]=32'h00000000;	data[347][9]=32'h3a1324e0;	data[347][10]=32'h38f7d209;	data[347][11]=32'h39aa60bc;	data[347][12]=32'h38f7d209;	data[347][13]=32'h00000000;	data[347][14]=32'h00000000;	data[347][15]=32'h00000000;	data[347][16]=32'h3a1324e0;
data[348][0]=32'h3b41cf43;	data[348][1]=32'h3f7ffa1a;	data[348][2]=32'h3c5b7ae5;	data[348][3]=32'h00000000;	data[348][4]=32'h39460e17;	data[348][5]=32'h37e27e0f;	data[348][6]=32'h39a9c25c;	data[348][7]=32'h00000000;	data[348][8]=32'h38e2587a;	data[348][9]=32'h38a9a8db;	data[348][10]=32'h00000000;	data[348][11]=32'h39460e17;	data[348][12]=32'h38a9a8db;	data[348][13]=32'h00000000;	data[348][14]=32'h37e27e0f;	data[348][15]=32'h00000000;	data[348][16]=32'h38a9a8db;
data[349][0]=32'h3b41ca3a;	data[349][1]=32'h3f7ffac2;	data[349][2]=32'h3c4aafbc;	data[349][3]=32'h00000000;	data[349][4]=32'h00000000;	data[349][5]=32'h00000000;	data[349][6]=32'h00000000;	data[349][7]=32'h3862e96f;	data[349][8]=32'h00000000;	data[349][9]=32'h00000000;	data[349][10]=32'h00000000;	data[349][11]=32'h00000000;	data[349][12]=32'h00000000;	data[349][13]=32'h00000000;	data[349][14]=32'h00000000;	data[349][15]=32'h3862e96f;	data[349][16]=32'h00000000;
data[350][0]=32'h3b705a71;	data[350][1]=32'h00000000;	data[350][2]=32'h3f6bce85;	data[350][3]=32'h394f90cc;	data[350][4]=32'h39c620e1;	data[350][5]=32'h390416d0;	data[350][6]=32'h00000000;	data[350][7]=32'h3896feb5;	data[350][8]=32'h38bcbe62;	data[350][9]=32'h39febc5e;	data[350][10]=32'h394f90cc;	data[350][11]=32'h39c620e1;	data[350][12]=32'h39754dca;	data[350][13]=32'h39a9d277;	data[350][14]=32'h390416d0;	data[350][15]=32'h3896feb5;	data[350][16]=32'h39febc5e;
data[351][0]=32'h3c6ad4f6;	data[351][1]=32'h00000000;	data[351][2]=32'h3f7c5586;	data[351][3]=32'h39daea9d;	data[351][4]=32'h3a007ec0;	data[351][5]=32'h39184b91;	data[351][6]=32'h00000000;	data[351][7]=32'h39e47002;	data[351][8]=32'h39b4d7b9;	data[351][9]=32'h39ab53ab;	data[351][10]=32'h39daea9d;	data[351][11]=32'h3a007ec0;	data[351][12]=32'h39184b91;	data[351][13]=32'h3a0ec580;	data[351][14]=32'h39184b91;	data[351][15]=32'h39e47002;	data[351][16]=32'h39ab53ab;
data[352][0]=32'h3d9c3bd6;	data[352][1]=32'h00000000;	data[352][2]=32'h3f7a656b;	data[352][3]=32'h3a2b3e32;	data[352][4]=32'h3a0d05e2;	data[352][5]=32'h39c97681;	data[352][6]=32'h39d388d4;	data[352][7]=32'h3a94954e;	data[352][8]=32'h3a355084;	data[352][9]=32'h3a5d9b26;	data[352][10]=32'h3a2b3e32;	data[352][11]=32'h3a0d05e2;	data[352][12]=32'h3a120f0c;	data[352][13]=32'h3a5388d4;	data[352][14]=32'h39c97681;	data[352][15]=32'h3a94954e;	data[352][16]=32'h3a5d9b26;
data[353][0]=32'h3b705a71;	data[353][1]=32'h00000000;	data[353][2]=32'h3f6bce85;	data[353][3]=32'h394f90cc;	data[353][4]=32'h39c620e1;	data[353][5]=32'h390416d0;	data[353][6]=32'h00000000;	data[353][7]=32'h3896feb5;	data[353][8]=32'h38bcbe62;	data[353][9]=32'h39febc5e;	data[353][10]=32'h394f90cc;	data[353][11]=32'h39c620e1;	data[353][12]=32'h39754dca;	data[353][13]=32'h39a9d277;	data[353][14]=32'h390416d0;	data[353][15]=32'h3896feb5;	data[353][16]=32'h39febc5e;
data[354][0]=32'h3b5e14f4;	data[354][1]=32'h00000000;	data[354][2]=32'h3f7f0260;	data[354][3]=32'h39907503;	data[354][4]=32'h3a61b76b;	data[354][5]=32'h379048b8;	data[354][6]=32'h00000000;	data[354][7]=32'h39349345;	data[354][8]=32'h38d8ad81;	data[354][9]=32'h396abea5;	data[354][10]=32'h39907503;	data[354][11]=32'h3a61b76b;	data[354][12]=32'h38fccfca;	data[354][13]=32'h38907e68;	data[354][14]=32'h379048b8;	data[354][15]=32'h39349345;	data[354][16]=32'h396abea5;
data[355][0]=32'h3c39c305;	data[355][1]=32'h3c9e16d7;	data[355][2]=32'h3f7fcb92;	data[355][3]=32'h397b8daa;	data[355][4]=32'h398fbe79;	data[355][5]=32'h38579654;	data[355][6]=32'h00000000;	data[355][7]=32'h39579e62;	data[355][8]=32'h380fdd58;	data[355][9]=32'h3933af1a;	data[355][10]=32'h397b8daa;	data[355][11]=32'h398fbe79;	data[355][12]=32'h39cea1e4;	data[355][13]=32'h3933af1a;	data[355][14]=32'h38579654;	data[355][15]=32'h39579e62;	data[355][16]=32'h3933af1a;
data[356][0]=32'h3c4cea29;	data[356][1]=32'h3c34e981;	data[356][2]=32'h3f7ff972;	data[356][3]=32'h39219df5;	data[356][4]=32'h38fb6816;	data[356][5]=32'h39339192;	data[356][6]=32'h396971c9;	data[356][7]=32'h380fdd58;	data[356][8]=32'h38b38426;	data[356][9]=32'h3998a2cf;	data[356][10]=32'h39219df5;	data[356][11]=32'h38fb6816;	data[356][12]=32'h397b6567;	data[356][13]=32'h38d77b7c;	data[356][14]=32'h39339192;	data[356][15]=32'h380fdd58;	data[356][16]=32'h3998a2cf;
data[357][0]=32'h3ecc9470;	data[357][1]=32'h00000000;	data[357][2]=32'h3f5bd513;	data[357][3]=32'h39200b4e;	data[357][4]=32'h39d20fad;	data[357][5]=32'h39960bc6;	data[357][6]=32'h39820a06;	data[357][7]=32'h39f0124c;	data[357][8]=32'h39dc108d;	data[357][9]=32'h39c80ecd;	data[357][10]=32'h39200b4e;	data[357][11]=32'h39d20fad;	data[357][12]=32'h395c108d;	data[357][13]=32'h39fa132c;	data[357][14]=32'h39960bc6;	data[357][15]=32'h39f0124c;	data[357][16]=32'h39c80ecd;
data[358][0]=32'h3e016c61;	data[358][1]=32'h00000000;	data[358][2]=32'h3f6b87be;	data[358][3]=32'h3905914f;	data[358][4]=32'h39abbb04;	data[358][5]=32'h3951e4ba;	data[358][6]=32'h3798ac34;	data[358][7]=32'h39abbb04;	data[358][8]=32'h39abbb04;	data[358][9]=32'h3a00cc99;	data[358][10]=32'h3905914f;	data[358][11]=32'h39abbb04;	data[358][12]=32'h398f1c12;	data[358][13]=32'h39abbb04;	data[358][14]=32'h3951e4ba;	data[358][15]=32'h39abbb04;	data[358][16]=32'h3a00cc99;
data[359][0]=32'h3c865732;	data[359][1]=32'h3cc3fe5d;	data[359][2]=32'h3f7fdd44;	data[359][3]=32'h398761b4;	data[359][4]=32'h392274b5;	data[359][5]=32'h381048b8;	data[359][6]=32'h381048b8;	data[359][7]=32'h39a274b5;	data[359][8]=32'h39589d66;	data[359][9]=32'h3a0be4a5;	data[359][10]=32'h398761b4;	data[359][11]=32'h392274b5;	data[359][12]=32'h39906797;	data[359][13]=32'h3934832a;	data[359][14]=32'h381048b8;	data[359][15]=32'h39a274b5;	data[359][16]=32'h3a0be4a5;
data[360][0]=32'h3d1ca07f;	data[360][1]=32'h3c217f41;	data[360][2]=32'h3f7ff972;	data[360][3]=32'h38d7b68b;	data[360][4]=32'h39c5bc37;	data[360][5]=32'h38b3b9d6;	data[360][6]=32'h38fba882;	data[360][7]=32'h39fba882;	data[360][8]=32'h3986d217;	data[360][9]=32'h39b3c1e4;	data[360][10]=32'h38d7b68b;	data[360][11]=32'h39c5bc37;	data[360][12]=32'h3998cb13;	data[360][13]=32'h3957b68b;	data[360][14]=32'h38b3b9d6;	data[360][15]=32'h39fba882;	data[360][16]=32'h39b3c1e4;
data[361][0]=32'h3c6c7c95;	data[361][1]=32'h00000000;	data[361][2]=32'h3f7705a7;	data[361][3]=32'h3a38a172;	data[361][4]=32'h399b7a44;	data[361][5]=32'h3a1b7a44;	data[361][6]=32'h399b7a44;	data[361][7]=32'h3a38a172;	data[361][8]=32'h39b8a21d;	data[361][9]=32'h39d5c89f;	data[361][10]=32'h3a38a172;	data[361][11]=32'h399b7a44;	data[361][12]=32'h391b7b9c;	data[361][13]=32'h3a5aa426;	data[361][14]=32'h3a1b7a44;	data[361][15]=32'h3a38a172;	data[361][16]=32'h39d5c89f;
data[362][0]=32'h3e33458d;	data[362][1]=32'h00000000;	data[362][2]=32'h3f605db7;	data[362][3]=32'h39a05bd6;	data[362][4]=32'h39be6be1;	data[362][5]=32'h38f08b18;	data[362][6]=32'h38a06ea0;	data[362][7]=32'h3a255e49;	data[362][8]=32'h39c8721f;	data[362][9]=32'h39f08869;	data[362][10]=32'h39a05bd6;	data[362][11]=32'h39be6be1;	data[362][12]=32'h395c7e9c;	data[362][13]=32'h3a074ce6;	data[362][14]=32'h38f08b18;	data[362][15]=32'h3a255e49;	data[362][16]=32'h39f08869;
data[363][0]=32'h3c216e0f;	data[363][1]=32'h00000000;	data[363][2]=32'h3f641893;	data[363][3]=32'h39f3d753;	data[363][4]=32'h3a146c5e;	data[363][5]=32'h39bed492;	data[363][6]=32'h39bed492;	data[363][7]=32'h3a09d27c;	data[363][8]=32'h387e9821;	data[363][9]=32'h397e6fdd;	data[363][10]=32'h39f3d753;	data[363][11]=32'h3a146c5e;	data[363][12]=32'h39693c19;	data[363][13]=32'h3a29a0ce;	data[363][14]=32'h39bed492;	data[363][15]=32'h3a09d27c;	data[363][16]=32'h397e6fdd;
data[364][0]=32'h3dd6e04c;	data[364][1]=32'h00000000;	data[364][2]=32'h3f750d06;	data[364][3]=32'h39f4582c;	data[364][4]=32'h3a3e96d4;	data[364][5]=32'h396a9103;	data[364][6]=32'h386a762b;	data[364][7]=32'h392fee1a;	data[364][8]=32'h39b9b3eb;	data[364][9]=32'h3a34d103;	data[364][10]=32'h39f4582c;	data[364][11]=32'h3a3e96d4;	data[364][12]=32'h39929b4e;	data[364][13]=32'h394379bd;	data[364][14]=32'h396a9103;	data[364][15]=32'h392fee1a;	data[364][16]=32'h3a34d103;
data[365][0]=32'h3d97e6f7;	data[365][1]=32'h00000000;	data[365][2]=32'h3f6cc2f8;	data[365][3]=32'h39a1f68a;	data[365][4]=32'h3a17d778;	data[365][5]=32'h394a7585;	data[365][6]=32'h395eb252;	data[365][7]=32'h39d493ec;	data[365][8]=32'h39f2f1d0;	data[365][9]=32'h3a0db865;	data[365][10]=32'h39a1f68a;	data[365][11]=32'h3a17d778;	data[365][12]=32'h3997d823;	data[365][13]=32'h39ac1649;	data[365][14]=32'h394a7585;	data[365][15]=32'h39d493ec;	data[365][16]=32'h3a0db865;
data[366][0]=32'h3d0e64b2;	data[366][1]=32'h3cf2580c;	data[366][2]=32'h3f7fc45d;	data[366][3]=32'h3999ca16;	data[366][4]=32'h38fd4b45;	data[366][5]=32'h38fd4b45;	data[366][6]=32'h3999ca16;	data[366][7]=32'h3910bed5;	data[366][8]=32'h3922d558;	data[366][9]=32'h39abe1f1;	data[366][10]=32'h3999ca16;	data[366][11]=32'h38fd4b45;	data[366][12]=32'h3934ee8a;	data[366][13]=32'h3922d558;	data[366][14]=32'h38fd4b45;	data[366][15]=32'h3910bed5;	data[366][16]=32'h39abe1f1;
data[367][0]=32'h3c33cc4b;	data[367][1]=32'h3c3ccaf7;	data[367][2]=32'h3f7ff62b;	data[367][3]=32'h388ed0e9;	data[367][4]=32'h00000000;	data[367][5]=32'h38d61927;	data[367][6]=32'h378e9b39;	data[367][7]=32'h388ed0e9;	data[367][8]=32'h39444061;	data[367][9]=32'h38f9c553;	data[367][10]=32'h388ed0e9;	data[367][11]=32'h00000000;	data[367][12]=32'h378e9b39;	data[367][13]=32'h39e7f095;	data[367][14]=32'h38d61927;	data[367][15]=32'h388ed0e9;	data[367][16]=32'h38f9c553;
data[368][0]=32'h3e4e8a72;	data[368][1]=32'h00000000;	data[368][2]=32'h3f73c6a8;	data[368][3]=32'h3a93a05b;	data[368][4]=32'h3a32435f;	data[368][5]=32'h3a2cb14e;	data[368][6]=32'h39c88ba0;	data[368][7]=32'h3a37d56f;	data[368][8]=32'h3a887c3b;	data[368][9]=32'h3a99326c;	data[368][10]=32'h3a93a05b;	data[368][11]=32'h3a32435f;	data[368][12]=32'h3a53afc0;	data[368][13]=32'h3ad6791e;	data[368][14]=32'h3a2cb14e;	data[368][15]=32'h3a37d56f;	data[368][16]=32'h3a99326c;
data[369][0]=32'h3d73a14d;	data[369][1]=32'h3d1bae47;	data[369][2]=32'h3f7dfaec;	data[369][3]=32'h39f0b0ad;	data[369][4]=32'h39d3ce9f;	data[369][5]=32'h3906c8b2;	data[369][6]=32'h38c084c0;	data[369][7]=32'h3986c8b2;	data[369][8]=32'h3986c8b2;	data[369][9]=32'h39ca2e62;	data[369][10]=32'h39f0b0ad;	data[369][11]=32'h39d3ce9f;	data[369][12]=32'h3953cd47;	data[369][13]=32'h3a0b997c;	data[369][14]=32'h3906c8b2;	data[369][15]=32'h3986c8b2;	data[369][16]=32'h39ca2e62;
data[370][0]=32'h3b953ec1;	data[370][1]=32'h00000000;	data[370][2]=32'h3f704578;	data[370][3]=32'h398494fb;	data[370][4]=32'h3a20fd91;	data[370][5]=32'h38979fc4;	data[370][6]=32'h00000000;	data[370][7]=32'h39763754;	data[370][8]=32'h39505771;	data[370][9]=32'h39c6de20;	data[370][10]=32'h398494fb;	data[370][11]=32'h3a20fd91;	data[370][12]=32'h38e34a12;	data[370][13]=32'h39ffb0a5;	data[370][14]=32'h38979fc4;	data[370][15]=32'h39763754;	data[370][16]=32'h39c6de20;
data[371][0]=32'h3cf676ea;	data[371][1]=32'h00000000;	data[371][2]=32'h3f769f6b;	data[371][3]=32'h39e2f025;	data[371][4]=32'h3a129091;	data[371][5]=32'h393d1f05;	data[371][6]=32'h3796feb5;	data[371][7]=32'h3975d961;	data[371][8]=32'h3975d961;	data[371][9]=32'h3a04614e;	data[371][10]=32'h39e2f025;	data[371][11]=32'h3a129091;	data[371][12]=32'h3975d961;	data[371][13]=32'h392a3471;	data[371][14]=32'h393d1f05;	data[371][15]=32'h3975d961;	data[371][16]=32'h3a04614e;
data[372][0]=32'h3df890d6;	data[372][1]=32'h3d324745;	data[372][2]=32'h3f7c3223;	data[372][3]=32'h3a0f6ff5;	data[372][4]=32'h3ae915d9;	data[372][5]=32'h3a001209;	data[372][6]=32'h3a42aa5f;	data[372][7]=32'h3ac01960;	data[372][8]=32'h39eba580;	data[372][9]=32'h3b0e2776;	data[372][10]=32'h3a0f6ff5;	data[372][11]=32'h3ae915d9;	data[372][12]=32'h3a148f44;	data[372][13]=32'h3b0a5050;	data[372][14]=32'h3a001209;	data[372][15]=32'h3ac01960;	data[372][16]=32'h3b0e2776;
data[373][0]=32'h3e8e7579;	data[373][1]=32'h00000000;	data[373][2]=32'h3f706c22;	data[373][3]=32'h389c7292;	data[373][4]=32'h3a8b687e;	data[373][5]=32'h3a0412ca;	data[373][6]=32'h381c7292;	data[373][7]=32'h39f49492;	data[373][8]=32'h3988f70a;	data[373][9]=32'h39573b10;	data[373][10]=32'h389c7292;	data[373][11]=32'h3a8b687e;	data[373][12]=32'h39fe5d13;	data[373][13]=32'h3a17a31f;	data[373][14]=32'h3a0412ca;	data[373][15]=32'h39f49492;	data[373][16]=32'h39573b10;
data[374][0]=32'h3ebe54b5;	data[374][1]=32'h00000000;	data[374][2]=32'h3f687dd4;	data[374][3]=32'h39d46ba8;	data[374][4]=32'h3a24a05e;	data[374][5]=32'h3a1f50be;	data[374][6]=32'h39d46ba8;	data[374][7]=32'h3a546ba8;	data[374][8]=32'h3969aa28;	data[374][9]=32'h3a6ef91d;	data[374][10]=32'h39d46ba8;	data[374][11]=32'h3a24a05e;	data[374][12]=32'h3a1f50be;	data[374][13]=32'h3a447d73;	data[374][14]=32'h3a1f50be;	data[374][15]=32'h3a546ba8;	data[374][16]=32'h3a6ef91d;
data[375][0]=32'h3e69e98e;	data[375][1]=32'h00000000;	data[375][2]=32'h3f742b95;	data[375][3]=32'h39e4b06e;	data[375][4]=32'h3987229f;	data[375][5]=32'h393b1b9f;	data[375][6]=32'h394fe6b3;	data[375][7]=32'h399bec5a;	data[375][8]=32'h3987229f;	data[375][9]=32'h39e4b06e;	data[375][10]=32'h39e4b06e;	data[375][11]=32'h3987229f;	data[375][12]=32'h39b0b76d;	data[375][13]=32'h3a1bed06;	data[375][14]=32'h393b1b9f;	data[375][15]=32'h399bec5a;	data[375][16]=32'h39e4b06e;
data[376][0]=32'h3c8904f7;	data[376][1]=32'h00000000;	data[376][2]=32'h3f7367a1;	data[376][3]=32'h3a231d26;	data[376][4]=32'h39efdf4b;	data[376][5]=32'h395316be;	data[376][6]=32'h39065544;	data[376][7]=32'h38e649cb;	data[376][8]=32'h393fe65f;	data[376][9]=32'h39c97e8f;	data[376][10]=32'h3a231d26;	data[376][11]=32'h39efdf4b;	data[376][12]=32'h39acb601;	data[376][13]=32'h39bfe65f;	data[376][14]=32'h395316be;	data[376][15]=32'h38e649cb;	data[376][16]=32'h39c97e8f;
data[377][0]=32'h3e6d3847;	data[377][1]=32'h00000000;	data[377][2]=32'h3f7421c0;	data[377][3]=32'h3a491dec;	data[377][4]=32'h3a33f235;	data[377][5]=32'h3a7374ac;	data[377][6]=32'h39de49a2;	data[377][7]=32'h3a96d671;	data[377][8]=32'h3a1ec67f;	data[377][9]=32'h3a1430a4;	data[377][10]=32'h3a491dec;	data[377][11]=32'h3a33f235;	data[377][12]=32'h39de49a2;	data[377][13]=32'h3a099b75;	data[377][14]=32'h3a7374ac;	data[377][15]=32'h3a96d671;	data[377][16]=32'h3a1430a4;
data[378][0]=32'h3e0e87d3;	data[378][1]=32'h00000000;	data[378][2]=32'h3f63ea0c;	data[378][3]=32'h39ac52af;	data[378][4]=32'h39192d0d;	data[378][5]=32'h00000000;	data[378][6]=32'h00000000;	data[378][7]=32'h3978e935;	data[378][8]=32'h39b5e580;	data[378][9]=32'h3a27889b;	data[378][10]=32'h39ac52af;	data[378][11]=32'h39192d0d;	data[378][12]=32'h3978e935;	data[378][13]=32'h39ac52af;	data[378][14]=32'h00000000;	data[378][15]=32'h3978e935;	data[378][16]=32'h3a27889b;
data[379][0]=32'h3d8cd749;	data[379][1]=32'h00000000;	data[379][2]=32'h3f6170f8;	data[379][3]=32'h39fc69c8;	data[379][4]=32'h39bfd644;	data[379][5]=32'h39b5bd3c;	data[379][6]=32'h39218b2b;	data[379][7]=32'h39de2006;	data[379][8]=32'h3a30b0b7;	data[379][9]=32'h39bfd644;	data[379][10]=32'h39fc69c8;	data[379][11]=32'h39bfd644;	data[379][12]=32'h395e1eaf;	data[379][13]=32'h3997737a;	data[379][14]=32'h39b5bd3c;	data[379][15]=32'h39de2006;	data[379][16]=32'h39bfd644;
data[380][0]=32'h3d6ba5a0;	data[380][1]=32'h3d8d3522;	data[380][2]=32'h3f7f1c97;	data[380][3]=32'h395fabf8;	data[380][4]=32'h3a027a18;	data[380][5]=32'h39d65aeb;	data[380][6]=32'h3a35bbe4;	data[380][7]=32'h39f24f68;	data[380][8]=32'h393a6516;	data[380][9]=32'h39fba1cc;	data[380][10]=32'h395fabf8;	data[380][11]=32'h3a027a18;	data[380][12]=32'h3982796c;	data[380][13]=32'h3a725014;	data[380][14]=32'h39d65aeb;	data[380][15]=32'h39f24f68;	data[380][16]=32'h39fba1cc;
data[381][0]=32'h3e9b4cc2;	data[381][1]=32'h00000000;	data[381][2]=32'h3f5f2b02;	data[381][3]=32'h391256da;	data[381][4]=32'h3a5b839f;	data[381][5]=32'h39bc280f;	data[381][6]=32'h391256da;	data[381][7]=32'h3a2c799b;	data[381][8]=32'h39925832;	data[381][9]=32'h399ccb27;	data[381][10]=32'h391256da;	data[381][11]=32'h3a5b839f;	data[381][12]=32'h39925832;	data[381][13]=32'h3a564978;	data[381][14]=32'h39bc280f;	data[381][15]=32'h3a2c799b;	data[381][16]=32'h399ccb27;
data[382][0]=32'h384d19fa;	data[382][1]=32'h00000000;	data[382][2]=32'h3f68ee8d;	data[382][3]=32'h39294ae8;	data[382][4]=32'h39967c84;	data[382][5]=32'h00000000;	data[382][6]=32'h00000000;	data[382][7]=32'h38bc1d52;	data[382][8]=32'h3961ba1a;	data[382][9]=32'h39eb21f7;	data[382][10]=32'h39294ae8;	data[382][11]=32'h39967c84;	data[382][12]=32'h397489d5;	data[382][13]=32'h39bc1aa3;	data[382][14]=32'h00000000;	data[382][15]=32'h38bc1d52;	data[382][16]=32'h39eb21f7;
data[383][0]=32'h3d5c5c57;	data[383][1]=32'h3d0257c9;	data[383][2]=32'h3f7faebc;	data[383][3]=32'h3970fe85;	data[383][4]=32'h399d91cc;	data[383][5]=32'h39b01bbc;	data[383][6]=32'h395e7495;	data[383][7]=32'h39d52e45;	data[383][8]=32'h398b07db;	data[383][9]=32'h398b07db;	data[383][10]=32'h3970fe85;	data[383][11]=32'h399d91cc;	data[383][12]=32'h398b07db;	data[383][13]=32'h394beaa5;	data[383][14]=32'h39b01bbc;	data[383][15]=32'h39d52e45;	data[383][16]=32'h398b07db;
data[384][0]=32'h3dad527e;	data[384][1]=32'h00000000;	data[384][2]=32'h3f6a1ff3;	data[384][3]=32'h394b011b;	data[384][4]=32'h3a03f497;	data[384][5]=32'h39739aed;	data[384][6]=32'h3936b432;	data[384][7]=32'h39cb011b;	data[384][8]=32'h39b6b432;	data[384][9]=32'h39226749;	data[384][10]=32'h394b011b;	data[384][11]=32'h3a03f497;	data[384][12]=32'h39a26749;	data[384][13]=32'h3a0907d1;	data[384][14]=32'h39739aed;	data[384][15]=32'h39cb011b;	data[384][16]=32'h39226749;
data[385][0]=32'h3d177425;	data[385][1]=32'h00000000;	data[385][2]=32'h3f7009d5;	data[385][3]=32'h398f343b;	data[385][4]=32'h38cc78ea;	data[385][5]=32'h39cc93c2;	data[385][6]=32'h38cc78ea;	data[385][7]=32'h39c2592b;	data[385][8]=32'h39381e95;	data[385][9]=32'h39ffb8b2;	data[385][10]=32'h398f343b;	data[385][11]=32'h38cc78ea;	data[385][12]=32'h398f343b;	data[385][13]=32'h3a04f9a4;	data[385][14]=32'h39cc93c2;	data[385][15]=32'h39c2592b;	data[385][16]=32'h39ffb8b2;
data[386][0]=32'h3b42b36e;	data[386][1]=32'h00000000;	data[386][2]=32'h3f794af5;	data[386][3]=32'h3950e058;	data[386][4]=32'h39f6db13;	data[386][5]=32'h39a16845;	data[386][6]=32'h3863c02e;	data[386][7]=32'h3a132a3f;	data[386][8]=32'h3963ddb5;	data[386][9]=32'h39aae6f4;	data[386][10]=32'h3950e058;	data[386][11]=32'h39f6db13;	data[386][12]=32'h3a04ec38;	data[386][13]=32'h3a17e996;	data[386][14]=32'h39a16845;	data[386][15]=32'h3a132a3f;	data[386][16]=32'h39aae6f4;
data[387][0]=32'h3d84894c;	data[387][1]=32'h3c50fa59;	data[387][2]=32'h3f7fa6df;	data[387][3]=32'h39f50aaf;	data[387][4]=32'h3a121516;	data[387][5]=32'h39750aaf;	data[387][6]=32'h39f50aaf;	data[387][7]=32'h3a16cbb4;	data[387][8]=32'h3a121516;	data[387][9]=32'h3a0d5e78;	data[387][10]=32'h39f50aaf;	data[387][11]=32'h3a121516;	data[387][12]=32'h39c5eb31;	data[387][13]=32'h39cf5716;	data[387][14]=32'h39750aaf;	data[387][15]=32'h3a16cbb4;	data[387][16]=32'h3a0d5e78;
data[388][0]=32'h3db9f98b;	data[388][1]=32'h00000000;	data[388][2]=32'h3f5efa83;	data[388][3]=32'h39f9fc5b;	data[388][4]=32'h39dd23b2;	data[388][5]=32'h39069b0f;	data[388][6]=32'h00000000;	data[388][7]=32'h3919d62a;	data[388][8]=32'h39869b0f;	data[388][9]=32'h39a373b8;	data[388][10]=32'h39f9fc5b;	data[388][11]=32'h39dd23b2;	data[388][12]=32'h392d1146;	data[388][13]=32'h39a373b8;	data[388][14]=32'h39069b0f;	data[388][15]=32'h3919d62a;	data[388][16]=32'h39a373b8;
data[389][0]=32'h3eadbb5a;	data[389][1]=32'h00000000;	data[389][2]=32'h3f4f0846;	data[389][3]=32'h3816feb5;	data[389][4]=32'h39b35e92;	data[389][5]=32'h39a07d64;	data[389][6]=32'h00000000;	data[389][7]=32'h3a381733;	data[389][8]=32'h39d92246;	data[389][9]=32'h39a9eea6;	data[389][10]=32'h3816feb5;	data[389][11]=32'h39b35e92;	data[389][12]=32'h3975735f;	data[389][13]=32'h38bcbe62;	data[389][14]=32'h39a07d64;	data[389][15]=32'h3a381733;	data[389][16]=32'h39a9eea6;
data[390][0]=32'h3e0f2a5a;	data[390][1]=32'h3d1ca9ef;	data[390][2]=32'h3f7e646f;	data[390][3]=32'h3a65c99e;	data[390][4]=32'h3a4d57b7;	data[390][5]=32'h39fe3b85;	data[390][6]=32'h3a8b57b7;	data[390][7]=32'h3a978efd;	data[390][8]=32'h39a63b13;	data[390][9]=32'h39cd57b7;	data[390][10]=32'h3a65c99e;	data[390][11]=32'h3a4d57b7;	data[390][12]=32'h39d71ee0;	data[390][13]=32'h3a9a0275;	data[390][14]=32'h39fe3b85;	data[390][15]=32'h3a978efd;	data[390][16]=32'h39cd57b7;
data[391][0]=32'h3cd2135e;	data[391][1]=32'h3d8d423e;	data[391][2]=32'h3f7f4e66;	data[391][3]=32'h39e77d27;	data[391][4]=32'h3994273f;	data[391][5]=32'h399d6988;	data[391][6]=32'h3901a2ad;	data[391][7]=32'h3994273f;	data[391][8]=32'h398ae4f6;	data[391][9]=32'h398ae4f6;	data[391][10]=32'h39e77d27;	data[391][11]=32'h3994273f;	data[391][12]=32'h3994273f;	data[391][13]=32'h3994273f;	data[391][14]=32'h399d6988;	data[391][15]=32'h3994273f;	data[391][16]=32'h398ae4f6;
data[392][0]=32'h3ccc7d1c;	data[392][1]=32'h3c74ba52;	data[392][2]=32'h3f7ff77b;	data[392][3]=32'h39973f21;	data[392][4]=32'h38f91ee5;	data[392][5]=32'h390e5acc;	data[392][6]=32'h38557d75;	data[392][7]=32'h398e5975;	data[392][8]=32'h39791c36;	data[392][9]=32'h38d58832;	data[392][10]=32'h39973f21;	data[392][11]=32'h38f91ee5;	data[392][12]=32'h388e6589;	data[392][13]=32'h388e6589;	data[392][14]=32'h390e5acc;	data[392][15]=32'h398e5975;	data[392][16]=32'h38d58832;
data[393][0]=32'h3b6aa01c;	data[393][1]=32'h00000000;	data[393][2]=32'h3f7128e1;	data[393][3]=32'h39b1c3dd;	data[393][4]=32'h39c47a18;	data[393][5]=32'h38e08ac5;	data[393][6]=32'h00000000;	data[393][7]=32'h39e08ac5;	data[393][8]=32'h3928696b;	data[393][9]=32'h398c5767;	data[393][10]=32'h39b1c3dd;	data[393][11]=32'h39c47a18;	data[393][12]=32'h39d73053;	data[393][13]=32'h39b1c3dd;	data[393][14]=32'h38e08ac5;	data[393][15]=32'h39e08ac5;	data[393][16]=32'h398c5767;
data[394][0]=32'h3cc56712;	data[394][1]=32'h3c195175;	data[394][2]=32'h3f7ffc11;	data[394][3]=32'h3984f197;	data[394][4]=32'h38b13598;	data[394][5]=32'h38b13598;	data[394][6]=32'h380dc479;	data[394][7]=32'h391f87c5;	data[394][8]=32'h388dc479;	data[394][9]=32'h38f827ef;	data[394][10]=32'h3984f197;	data[394][11]=32'h38b13598;	data[394][12]=32'h38d4b6d1;	data[394][13]=32'h39314304;	data[394][14]=32'h38b13598;	data[394][15]=32'h391f87c5;	data[394][16]=32'h38f827ef;
data[395][0]=32'h3c7f151e;	data[395][1]=32'h3c837718;	data[395][2]=32'h3f7ff4dc;	data[395][3]=32'h38b2e317;	data[395][4]=32'h39568f43;	data[395][5]=32'h380f0699;	data[395][6]=32'h38fa50e9;	data[395][7]=32'h39df7fad;	data[395][8]=32'h39a0eb72;	data[395][9]=32'h3920ea1b;	data[395][10]=32'h38b2e317;	data[395][11]=32'h39568f43;	data[395][12]=32'h38fa50e9;	data[395][13]=32'h39568f43;	data[395][14]=32'h380f0699;	data[395][15]=32'h39df7fad;	data[395][16]=32'h3920ea1b;
data[396][0]=32'h3db09635;	data[396][1]=32'h00000000;	data[396][2]=32'h3f7ef1fe;	data[396][3]=32'h3a147873;	data[396][4]=32'h3a22d603;	data[396][5]=32'h39861a36;	data[396][6]=32'h38e5e3ca;	data[396][7]=32'h3a7dd583;	data[396][8]=32'h39d2bb79;	data[396][9]=32'h3a194287;	data[396][10]=32'h3a147873;	data[396][11]=32'h3a22d603;	data[396][12]=32'h39861a36;	data[396][13]=32'h3a7dd583;	data[396][14]=32'h39861a36;	data[396][15]=32'h3a7dd583;	data[396][16]=32'h3a194287;
data[397][0]=32'h3c367c28;	data[397][1]=32'h3ca0125a;	data[397][2]=32'h3f7feda6;	data[397][3]=32'h38572af5;	data[397][4]=32'h38d7406e;	data[397][5]=32'h38b34e77;	data[397][6]=32'h378f71f8;	data[397][7]=32'h38b34e77;	data[397][8]=32'h38b34e77;	data[397][9]=32'h38b34e77;	data[397][10]=32'h38572af5;	data[397][11]=32'h38d7406e;	data[397][12]=32'h38fb224b;	data[397][13]=32'h38572af5;	data[397][14]=32'h38b34e77;	data[397][15]=32'h38b34e77;	data[397][16]=32'h38b34e77;
data[398][0]=32'h3c4065b6;	data[398][1]=32'h00000000;	data[398][2]=32'h3f725aee;	data[398][3]=32'h39e38520;	data[398][4]=32'h3a7ff670;	data[398][5]=32'h3817d574;	data[398][6]=32'h393d9a80;	data[398][7]=32'h3904b7e0;	data[398][8]=32'h39a12930;	data[398][9]=32'h39da0a78;	data[398][10]=32'h39e38520;	data[398][11]=32'h3a7ff670;	data[398][12]=32'h39e38520;	data[398][13]=32'h39ed0120;	data[398][14]=32'h3817d574;	data[398][15]=32'h3904b7e0;	data[398][16]=32'h39da0a78;
data[399][0]=32'h3b257c26;	data[399][1]=32'h00000000;	data[399][2]=32'h3f6ca57a;	data[399][3]=32'h397e1f55;	data[399][4]=32'h396a9103;	data[399][5]=32'h392fee1a;	data[399][6]=32'h379c0732;	data[399][7]=32'h3988d57c;	data[399][8]=32'h38ea9103;	data[399][9]=32'h397e1f55;	data[399][10]=32'h397e1f55;	data[399][11]=32'h396a9103;	data[399][12]=32'h39a626f1;	data[399][13]=32'h39a626f1;	data[399][14]=32'h392fee1a;	data[399][15]=32'h3988d57c;	data[399][16]=32'h397e1f55;
data[400][0]=32'h3d25bb7b;	data[400][1]=32'h3d109071;	data[400][2]=32'h3f7fce31;	data[400][3]=32'h399397a2;	data[400][4]=32'h3a1834c0;	data[400][5]=32'h3a01252f;	data[400][6]=32'h399cd1dd;	data[400][7]=32'h3a1cd1dd;	data[400][8]=32'h3a0efb30;	data[400][9]=32'h3a216e4f;	data[400][10]=32'h399397a2;	data[400][11]=32'h3a1834c0;	data[400][12]=32'h391398fa;	data[400][13]=32'h39c1b81c;	data[400][14]=32'h3a01252f;	data[400][15]=32'h3a1cd1dd;	data[400][16]=32'h3a216e4f;
data[401][0]=32'h3d6a5f85;	data[401][1]=32'h00000000;	data[401][2]=32'h3f765f31;	data[401][3]=32'h393dd83d;	data[401][4]=32'h3963d04a;	data[401][5]=32'h393dd83d;	data[401][6]=32'h3797d574;	data[401][7]=32'h3904e582;	data[401][8]=32'h3897d574;	data[401][9]=32'h3a261e37;	data[401][10]=32'h393dd83d;	data[401][11]=32'h3963d04a;	data[401][12]=32'h3963d04a;	data[401][13]=32'h39bdd995;	data[401][14]=32'h393dd83d;	data[401][15]=32'h3904e582;	data[401][16]=32'h3a261e37;
data[402][0]=32'h3d91ec0b;	data[402][1]=32'h00000000;	data[402][2]=32'h3f73f9c6;	data[402][3]=32'h3a095452;	data[402][4]=32'h39fe50fe;	data[402][5]=32'h3922c28d;	data[402][6]=32'h39c1475e;	data[402][7]=32'h3a2cef0c;	data[402][8]=32'h39843f14;	data[402][9]=32'h3a41475e;	data[402][10]=32'h3a095452;	data[402][11]=32'h39fe50fe;	data[402][12]=32'h38f42683;	data[402][13]=32'h3a5089c6;	data[402][14]=32'h3922c28d;	data[402][15]=32'h3a2cef0c;	data[402][16]=32'h3a41475e;
data[403][0]=32'h3b30aa57;	data[403][1]=32'h00000000;	data[403][2]=32'h3f712253;	data[403][3]=32'h39748477;	data[403][4]=32'h3916787d;	data[403][5]=32'h3916787d;	data[403][6]=32'h00000000;	data[403][7]=32'h3961b4bb;	data[403][8]=32'h38bc1d52;	data[403][9]=32'h38e1b76b;	data[403][10]=32'h39748477;	data[403][11]=32'h3916787d;	data[403][12]=32'h00000000;	data[403][13]=32'h39f48477;	data[403][14]=32'h3916787d;	data[403][15]=32'h3961b4bb;	data[403][16]=32'h38e1b76b;
data[404][0]=32'h3c916ebd;	data[404][1]=32'h00000000;	data[404][2]=32'h3f64ce1c;	data[404][3]=32'h39d39b9e;	data[404][4]=32'h39dd3a83;	data[404][5]=32'h39a383d3;	data[404][6]=32'h3819ee53;	data[404][7]=32'h3999e646;	data[404][8]=32'h39904760;	data[404][9]=32'h39f076f6;	data[404][10]=32'h39d39b9e;	data[404][11]=32'h39dd3a83;	data[404][12]=32'h392d2161;	data[404][13]=32'h3999e646;	data[404][14]=32'h39a383d3;	data[404][15]=32'h3999e646;	data[404][16]=32'h39f076f6;
data[405][0]=32'h3db99d45;	data[405][1]=32'h00000000;	data[405][2]=32'h3f721577;	data[405][3]=32'h39e45681;	data[405][4]=32'h3a86ecef;	data[405][5]=32'h3a2b40e1;	data[405][6]=32'h39c53350;	data[405][7]=32'h3aa37916;	data[405][8]=32'h3a73e81a;	data[405][9]=32'h3a0c1db0;	data[405][10]=32'h39e45681;	data[405][11]=32'h3a86ecef;	data[405][12]=32'h3a3071a2;	data[405][13]=32'h3a2b40e1;	data[405][14]=32'h3a2b40e1;	data[405][15]=32'h3aa37916;	data[405][16]=32'h3a0c1db0;
data[406][0]=32'h3b705a71;	data[406][1]=32'h00000000;	data[406][2]=32'h3f6bce85;	data[406][3]=32'h394f90cc;	data[406][4]=32'h39c620e1;	data[406][5]=32'h390416d0;	data[406][6]=32'h00000000;	data[406][7]=32'h3896feb5;	data[406][8]=32'h38bcbe62;	data[406][9]=32'h39febc5e;	data[406][10]=32'h394f90cc;	data[406][11]=32'h39c620e1;	data[406][12]=32'h39754dca;	data[406][13]=32'h39a9d277;	data[406][14]=32'h390416d0;	data[406][15]=32'h3896feb5;	data[406][16]=32'h39febc5e;
data[407][0]=32'h3da9f623;	data[407][1]=32'h00000000;	data[407][2]=32'h3f752e73;	data[407][3]=32'h3a0c205f;	data[407][4]=32'h3a2b443c;	data[407][5]=32'h3a6ebc0b;	data[407][6]=32'h3a01bf88;	data[407][7]=32'h3a4f982e;	data[407][8]=32'h3a791d8e;	data[407][9]=32'h3aa37c71;	data[407][10]=32'h3a0c205f;	data[407][11]=32'h3a2b443c;	data[407][12]=32'h3a8c210b;	data[407][13]=32'h3a73eccc;	data[407][14]=32'h3a6ebc0b;	data[407][15]=32'h3a4f982e;	data[407][16]=32'h3aa37c71;
data[408][0]=32'h3d067f0b;	data[408][1]=32'h3cc0ebee;	data[408][2]=32'h3f7feb07;	data[408][3]=32'h395547c6;	data[408][4]=32'h388e2fd9;	data[408][5]=32'h39670dc1;	data[408][6]=32'h00000000;	data[408][7]=32'h390e2fd9;	data[408][8]=32'h3931bbcf;	data[408][9]=32'h394381ca;	data[408][10]=32'h395547c6;	data[408][11]=32'h388e2fd9;	data[408][12]=32'h390e2fd9;	data[408][13]=32'h3931bbcf;	data[408][14]=32'h39670dc1;	data[408][15]=32'h390e2fd9;	data[408][16]=32'h394381ca;
data[409][0]=32'h3deaf252;	data[409][1]=32'h00000000;	data[409][2]=32'h3f7631f9;	data[409][3]=32'h39ebe89c;	data[409][4]=32'h39ebe89c;	data[409][5]=32'h379cddf2;	data[409][6]=32'h00000000;	data[409][7]=32'h39a719e0;	data[409][8]=32'h39e21407;	data[409][9]=32'h3a8e8717;	data[409][10]=32'h39ebe89c;	data[409][11]=32'h39ebe89c;	data[409][12]=32'h39ebe89c;	data[409][13]=32'h38ebe89c;	data[409][14]=32'h379cddf2;	data[409][15]=32'h39a719e0;	data[409][16]=32'h3a8e8717;
data[410][0]=32'h3dfaebc4;	data[410][1]=32'h00000000;	data[410][2]=32'h3f74b09f;	data[410][3]=32'h39cb2c0e;	data[410][4]=32'h391acd20;	data[410][5]=32'h392e25c3;	data[410][6]=32'h00000000;	data[410][7]=32'h391acd20;	data[410][8]=32'h39c17fbd;	data[410][9]=32'h3a3ca8e8;	data[410][10]=32'h39cb2c0e;	data[410][11]=32'h391acd20;	data[410][12]=32'h39911f78;	data[410][13]=32'h3a2e25c3;	data[410][14]=32'h392e25c3;	data[410][15]=32'h391acd20;	data[410][16]=32'h3a3ca8e8;
data[411][0]=32'h3cc3f812;	data[411][1]=32'h00000000;	data[411][2]=32'h3f5b81d8;	data[411][3]=32'h3a1f9485;	data[411][4]=32'h39a98e03;	data[411][5]=32'h390ba0de;	data[411][6]=32'h379f6230;	data[411][7]=32'h399f93da;	data[411][8]=32'h3a427cbd;	data[411][9]=32'h3a6a6209;	data[411][10]=32'h3a1f9485;	data[411][11]=32'h39a98e03;	data[411][12]=32'h398ba235;	data[411][13]=32'h39b386d6;	data[411][14]=32'h390ba0de;	data[411][15]=32'h399f93da;	data[411][16]=32'h3a6a6209;
data[412][0]=32'h3cd7f51f;	data[412][1]=32'h3cb24a6b;	data[412][2]=32'h3f7fe133;	data[412][3]=32'h39335e92;	data[412][4]=32'h38fb1cec;	data[412][5]=32'h38fb1cec;	data[412][6]=32'h38b34e77;	data[412][7]=32'h39454f80;	data[412][8]=32'h378f71f8;	data[412][9]=32'h398686ed;	data[412][10]=32'h39335e92;	data[412][11]=32'h38fb1cec;	data[412][12]=32'h390f7f64;	data[412][13]=32'h39aa661b;	data[412][14]=32'h38fb1cec;	data[412][15]=32'h39454f80;	data[412][16]=32'h398686ed;
data[413][0]=32'h3d6acd9f;	data[413][1]=32'h00000000;	data[413][2]=32'h3f78dae4;	data[413][3]=32'h3a2d22b8;	data[413][4]=32'h3a19e646;	data[413][5]=32'h392d2410;	data[413][6]=32'h3966d811;	data[413][7]=32'h3a31f22b;	data[413][8]=32'h39a3852b;	data[413][9]=32'h39ad22b8;	data[413][10]=32'h3a2d22b8;	data[413][11]=32'h3a19e646;	data[413][12]=32'h3986a9d3;	data[413][13]=32'h392d2410;	data[413][14]=32'h392d2410;	data[413][15]=32'h3a31f22b;	data[413][16]=32'h39ad22b8;
data[414][0]=32'h3ccddb55;	data[414][1]=32'h3cbd2d88;	data[414][2]=32'h3f7fe5c9;	data[414][3]=32'h380f0699;	data[414][4]=32'h3944a104;	data[414][5]=32'h00000000;	data[414][6]=32'h380f0699;	data[414][7]=32'h397a40ce;	data[414][8]=32'h388f0699;	data[414][9]=32'h38fa40ce;	data[414][10]=32'h380f0699;	data[414][11]=32'h3944a104;	data[414][12]=32'h38565435;	data[414][13]=32'h3997f1a4;	data[414][14]=32'h00000000;	data[414][15]=32'h397a40ce;	data[414][16]=32'h38fa40ce;
data[415][0]=32'h3ddd0fa6;	data[415][1]=32'h00000000;	data[415][2]=32'h3f68d25f;	data[415][3]=32'h39d9f7ae;	data[415][4]=32'h3a6457d9;	data[415][5]=32'h393ad325;	data[415][6]=32'h393ad325;	data[415][7]=32'h39bad325;	data[415][8]=32'h39645930;	data[415][9]=32'h3a2b4239;	data[415][10]=32'h39d9f7ae;	data[415][11]=32'h3a6457d9;	data[415][12]=32'h3a20e0b6;	data[415][13]=32'h39b072fa;	data[415][14]=32'h393ad325;	data[415][15]=32'h39bad325;	data[415][16]=32'h3a2b4239;
data[416][0]=32'h3c93d966;	data[416][1]=32'h3c58cf3a;	data[416][2]=32'h3f7ff823;	data[416][3]=32'h38b1a0f7;	data[416][4]=32'h390e27cb;	data[416][5]=32'h38f8c8ff;	data[416][6]=32'h38551216;	data[416][7]=32'h39670304;	data[416][8]=32'h38b1a0f7;	data[416][9]=32'h388e2fd9;	data[416][10]=32'h38b1a0f7;	data[416][11]=32'h390e27cb;	data[416][12]=32'h38b1a0f7;	data[416][13]=32'h39553d09;	data[416][14]=32'h38f8c8ff;	data[416][15]=32'h39670304;	data[416][16]=32'h388e2fd9;
data[417][0]=32'h3d51dde3;	data[417][1]=32'h3c170a73;	data[417][2]=32'h3f7fee4e;	data[417][3]=32'h39483711;	data[417][4]=32'h39a3cefd;	data[417][5]=32'h3923cefd;	data[417][6]=32'h39d14fbe;	data[417][7]=32'h39a3cefd;	data[417][8]=32'h396c9c76;	data[417][9]=32'h39c835b9;	data[417][10]=32'h39483711;	data[417][11]=32'h39a3cefd;	data[417][12]=32'h39483711;	data[417][13]=32'h39e383c8;	data[417][14]=32'h3923cefd;	data[417][15]=32'h39a3cefd;	data[417][16]=32'h39c835b9;
data[418][0]=32'h3c5cb9aa;	data[418][1]=32'h3cae9036;	data[418][2]=32'h3f7fdf3b;	data[418][3]=32'h390ff023;	data[418][4]=32'h39cee907;	data[418][5]=32'h38d7e6dc;	data[418][6]=32'h385801b4;	data[418][7]=32'h38d7e6dc;	data[418][8]=32'h38fbe391;	data[418][9]=32'h3957e6dc;	data[418][10]=32'h390ff023;	data[418][11]=32'h39cee907;	data[418][12]=32'h380fdd58;	data[418][13]=32'h390ff023;	data[418][14]=32'h38d7e6dc;	data[418][15]=32'h38d7e6dc;	data[418][16]=32'h3957e6dc;
data[419][0]=32'h3c2d2136;	data[419][1]=32'h3ce5d399;	data[419][2]=32'h3f7fb891;	data[419][3]=32'h381048b8;	data[419][4]=32'h396a88f5;	data[419][5]=32'h389048b8;	data[419][6]=32'h00000000;	data[419][7]=32'h39467418;	data[419][8]=32'h38b45ae6;	data[419][9]=32'h39105375;	data[419][10]=32'h381048b8;	data[419][11]=32'h396a88f5;	data[419][12]=32'h39105375;	data[419][13]=32'h39874ee9;	data[419][14]=32'h389048b8;	data[419][15]=32'h39467418;	data[419][16]=32'h39105375;
data[420][0]=32'h3d36deb9;	data[420][1]=32'h3d1dfdac;	data[420][2]=32'h3f7f6556;	data[420][3]=32'h3a05751f;	data[420][4]=32'h3a0a3929;	data[420][5]=32'h3a51b7c3;	data[420][6]=32'h39ee50ab;	data[420][7]=32'h3a13c13d;	data[420][8]=32'h39b51edb;	data[420][9]=32'h3a436ba5;	data[420][10]=32'h3a05751f;	data[420][11]=32'h3a0a3929;	data[420][12]=32'h3a3ea6ef;	data[420][13]=32'h3a8c99d7;	data[420][14]=32'h3a51b7c3;	data[420][15]=32'h3a13c13d;	data[420][16]=32'h3a436ba5;
data[421][0]=32'h3e93b3a7;	data[421][1]=32'h00000000;	data[421][2]=32'h3f66f7e4;	data[421][3]=32'h3a162749;	data[421][4]=32'h39b654e6;	data[421][5]=32'h39a0e0b6;	data[421][6]=32'h392b9976;	data[421][7]=32'h3a10ca3d;	data[421][8]=32'h3a0b6ddd;	data[421][9]=32'h3a0b6ddd;	data[421][10]=32'h3a162749;	data[421][11]=32'h39b654e6;	data[421][12]=32'h39c10da7;	data[421][13]=32'h3a30f7da;	data[421][14]=32'h39a0e0b6;	data[421][15]=32'h3a10ca3d;	data[421][16]=32'h3a0b6ddd;
data[422][0]=32'h3d083559;	data[422][1]=32'h3cd436b9;	data[422][2]=32'h3f7fe7c0;	data[422][3]=32'h39217302;	data[422][4]=32'h38572af5;	data[422][5]=32'h393363f0;	data[422][6]=32'h39aa6b79;	data[422][7]=32'h3957431d;	data[422][8]=32'h39217302;	data[422][9]=32'h38fb224b;	data[422][10]=32'h39217302;	data[422][11]=32'h38572af5;	data[422][12]=32'h380f71f8;	data[422][13]=32'h393363f0;	data[422][14]=32'h393363f0;	data[422][15]=32'h3957431d;	data[422][16]=32'h38fb224b;
data[423][0]=32'h3cb20fb2;	data[423][1]=32'h3c719d67;	data[423][2]=32'h3f7ff4dc;	data[423][3]=32'h390ec37d;	data[423][4]=32'h388ed0e9;	data[423][5]=32'h38b277b7;	data[423][6]=32'h388ed0e9;	data[423][7]=32'h38b277b7;	data[423][8]=32'h39209c42;	data[423][9]=32'h39a09c42;	data[423][10]=32'h390ec37d;	data[423][11]=32'h388ed0e9;	data[423][12]=32'h380e9b39;	data[423][13]=32'h390ec37d;	data[423][14]=32'h38b277b7;	data[423][15]=32'h38b277b7;	data[423][16]=32'h39a09c42;
data[424][0]=32'h3e1f1412;	data[424][1]=32'h00000000;	data[424][2]=32'h3f6b61bb;	data[424][3]=32'h3a32928f;	data[424][4]=32'h3a09c1b5;	data[424][5]=32'h3a09c1b5;	data[424][6]=32'h3823288f;	data[424][7]=32'h3a0edba6;	data[424][8]=32'h39990f86;	data[424][9]=32'h39e07eb0;	data[424][10]=32'h3a32928f;	data[424][11]=32'h3a09c1b5;	data[424][12]=32'h39607d59;	data[424][13]=32'h39ff1a52;	data[424][14]=32'h3a09c1b5;	data[424][15]=32'h3a0edba6;	data[424][16]=32'h39e07eb0;
data[425][0]=32'h3dae79ab;	data[425][1]=32'h00000000;	data[425][2]=32'h3f7557bc;	data[425][3]=32'h38e15c26;	data[425][4]=32'h39163d6f;	data[425][5]=32'h398cd998;	data[425][6]=32'h398cd998;	data[425][7]=32'h39f4252b;	data[425][8]=32'h379627f5;	data[425][9]=32'h398375c1;	data[425][10]=32'h38e15c26;	data[425][11]=32'h39163d6f;	data[425][12]=32'h39163d6f;	data[425][13]=32'h3a4e9524;	data[425][14]=32'h398cd998;	data[425][15]=32'h39f4252b;	data[425][16]=32'h398375c1;
data[426][0]=32'h3a13f037;	data[426][1]=32'h00000000;	data[426][2]=32'h3f54ab60;	data[426][3]=32'h379c0732;	data[426][4]=32'h3a209638;	data[426][5]=32'h00000000;	data[426][6]=32'h392f2f83;	data[426][7]=32'h39561e85;	data[426][8]=32'h389bd182;	data[426][9]=32'h399bb802;	data[426][10]=32'h379c0732;	data[426][11]=32'h3a209638;	data[426][12]=32'h38e994af;	data[426][13]=32'h392f2f83;	data[426][14]=32'h00000000;	data[426][15]=32'h39561e85;	data[426][16]=32'h399bb802;
data[427][0]=32'h3dea0126;	data[427][1]=32'h3ddfd8ae;	data[427][2]=32'h3f7d8cd2;	data[427][3]=32'h39990778;	data[427][4]=32'h3a0f76ab;	data[427][5]=32'h39ef1b56;	data[427][6]=32'h39190778;	data[427][7]=32'h39d2699a;	data[427][8]=32'h398f75ff;	data[427][9]=32'h398f75ff;	data[427][10]=32'h39990778;	data[427][11]=32'h3a0f76ab;	data[427][12]=32'h39990778;	data[427][13]=32'h3a143ebc;	data[427][14]=32'h39ef1b56;	data[427][15]=32'h39d2699a;	data[427][16]=32'h398f75ff;
data[428][0]=32'h3bd3be59;	data[428][1]=32'h3bc90314;	data[428][2]=32'h3f7ffe09;	data[428][3]=32'h388d236a;	data[428][4]=32'h391ebe72;	data[428][5]=32'h38d3aa62;	data[428][6]=32'h00000000;	data[428][7]=32'h38f6f08d;	data[428][8]=32'h388d236a;	data[428][9]=32'h38b05ed8;	data[428][10]=32'h388d236a;	data[428][11]=32'h391ebe72;	data[428][12]=32'h38b05ed8;	data[428][13]=32'h398449d1;	data[428][14]=32'h38d3aa62;	data[428][15]=32'h38f6f08d;	data[428][16]=32'h38b05ed8;
data[429][0]=32'h3d9d859d;	data[429][1]=32'h3d3a9b07;	data[429][2]=32'h3f7e1da8;	data[429][3]=32'h3a3b1844;	data[429][4]=32'h39efddf4;	data[429][5]=32'h389982f3;	data[429][6]=32'h389982f3;	data[429][7]=32'h398feac4;	data[429][8]=32'h3a4e48a3;	data[429][9]=32'h3a57e0d2;	data[429][10]=32'h3a3b1844;	data[429][11]=32'h39efddf4;	data[429][12]=32'h3966446d;	data[429][13]=32'h3a0b1f58;	data[429][14]=32'h389982f3;	data[429][15]=32'h398feac4;	data[429][16]=32'h3a57e0d2;
end


initial begin
    start_fix_conv = 0;
    reset = 1;
    @(posedge clk);
    reset = 0;
    for(int i=0; i<430; i++) begin //LBP_161, LBP_156, LBP_137, LBP_136, LBP_132, LBP_128, LBP_125, LBP_43, LBP_38, LBP_32, LBP_25, LBP_19, LBP_14, LBP_7
    b_bin208  = data[i][0];
    a_bin199  = data[i][1];
    a_bin198  = data[i][2];
    LBP_161   = data[i][3]; 
    LBP_156   = data[i][4];
    LBP_137   = data[i][5];	
    LBP_136   = data[i][6];
    LBP_132   = data[i][7];	
    LBP_128   = data[i][8];		
    LBP_125   = data[i][9];		
    LBP_43    = data[i][10];		
    LBP_38    = data[i][11];
    LBP_32    = data[i][12];		
    LBP_25    = data[i][13];		
    LBP_19    = data[i][14];	
    LBP_14    = data[i][15];		
    LBP_7     = data[i][16];
    start_fix_conv = 1;
    @(posedge clk);
    start_fix_conv = 0;
    repeat(35000) @(posedge clk);
    end
    $finish();
end
/*
initial begin
   clk = 0;
   reset = 1;
   # 10;
   reset = 0;
   start_fix_conv = 1;
   #10;
   start_fix_conv = 0;
   //both positive


   b_bin208 = 0.17507	;
   a_bin199 = 0	        ;
   a_bin198 = 0.87643	;
   LBP_161  = 0.00030586;		
   LBP_156  = 0.0003632	;
   LBP_137  = 0.0001147	;	
   LBP_136  = 7.65E-05	;	
   LBP_132  = 0.00063083;	
   LBP_128  = 0.00038232;		
   LBP_125  = 0.00045878;		
   LBP_43   = 0.00030586;		
   LBP_38   = 0.0003632	;
   LBP_32   = 0.00021028;		
   LBP_25   = 0.00051613;		
   LBP_19   = 0.0001147	;	
   LBP_14   = 0.00063083;		
   LBP_7    = 0.00045878;
/*
    LBP_166 = 32'h3b97a5a4;
    LBP_162 = 32'h3b8a48c4;
    LBP_161 = 32'h3b15a518;
    LBP_156 = 32'h3b41bb21; 
    LBP_150 = 32'h3b1c52b1;
    LBP_143 = 32'h3b3f104c;
    LBP_137 = 32'h3b1da8f3;
    LBP_136 = 32'h3af88334;
    LBP_132 = 32'h3b4dc1bf;
    LBP_131 = 32'h3ab5b482;
    LBP_125 = 32'h3b345fee;
    LBP_84  = 32'h3b0e3187;
    LBP_66  = 32'h3b11deba;
    LBP_43  = 32'h3b15a518;
    LBP_38  = 32'h3b41bb21;
    LBP_32  = 32'h3b1c52b1;
    LBP_25  = 32'h3b3f104c;
    LBP_19  = 32'h3b1da8f3;
    LBP_18  = 32'h3af88334;
    LBP_14  = 32'h3b4dc1bf;
    LBP_10  = 32'h3b0d9f90;
    LBP_7   = 32'h3b345fee;
    #100;
    


b_bin208 = 32'h3992ccf7;
a_bin199 = 32'h00000000; 
a_bin198 = 32'h3f5e65bf; //0.86874
LBP_161  = 32'h39e41365; //0.00043502
LBP_156  = 32'h3a2dc5cb; //0.00066289
LBP_137  = 32'h3a53c895; //0.00080789
LBP_136  = 32'h3a07c257; //0.00051788
LBP_132  = 32'h3abe1148; //0.0014501
LBP_128  = 32'h3a07c257; //0.00051788
LBP_125  = 32'h3a9ac513; //0.0011808
LBP_43   = 32'h39e41365; //0.00043502
LBP_38   = 32'h3a2dc5cb; //0.00066289
LBP_32   = 32'h398253d8; //0.00024858
LBP_25   = 32'h3ad112ad; //0.0015951
LBP_19   = 32'h3a53c895; //0.00080789
LBP_14   = 32'h3abe1148; //0.0014501
LBP_7    = 32'h3a9ac513; //0.0011808

end
*/
Fix_NN uut(.*);

endmodule

